magic
tech sky130A
magscale 1 2
timestamp 1700276902
<< error_p >>
rect 53968 3350 54640 4550
rect 56240 3350 57840 4550
rect 57900 3350 59500 4550
rect 61100 3350 62700 4550
rect 54700 1610 56300 2810
rect 54700 0 56300 1200
rect 56360 0 56547 1200
<< nwell >>
rect -4920 3280 67560 5050
rect -4920 3200 32120 3280
rect -4920 1770 27450 3200
<< nmos >>
rect 33780 1610 35380 2810
rect 38640 1610 40240 2810
rect 41840 1610 43440 2810
rect 45040 1610 46640 2810
rect 48240 1610 49840 2810
rect 53100 1610 54700 2810
rect 56300 1610 57900 2810
rect -3200 0 -1600 1200
rect 0 0 1600 1200
rect 4860 0 6460 1200
rect 8060 0 9660 1200
rect 12920 0 14520 1200
rect 16120 0 17720 1200
rect 20980 0 22580 1200
rect 24180 0 25780 1200
rect 27380 0 28980 1200
rect 30580 0 32180 1200
rect 33780 0 35380 1200
rect 36980 0 38580 1200
rect 41840 0 43440 1200
rect 45040 0 46640 1200
rect 49900 0 51500 1200
rect 53100 0 54700 1200
rect 57960 0 59560 1200
rect 61160 0 62760 1200
<< pmos >>
rect -1660 3350 -60 4550
rect 1540 3350 3140 4550
rect 6400 3350 8000 4550
rect 9600 3350 11200 4550
rect 14460 3350 16060 4550
rect 17660 3350 19260 4550
rect 22520 3350 24120 4550
rect 25720 3350 27320 4550
rect 28920 3350 30520 4550
rect 32120 3350 33720 4550
rect 35320 3350 36920 4550
rect 38520 3350 40120 4550
rect 43380 3350 44980 4550
rect 46580 3350 48180 4550
rect 51440 3350 53040 4550
rect 54640 3350 56240 4550
rect 59500 3350 61100 4550
rect 62700 3350 64300 4550
rect -1660 1810 -60 3010
rect 1540 1810 3140 3010
rect 6400 1810 8000 3010
rect 11260 1810 12860 3010
rect 14460 1810 16060 3010
rect 19320 1810 20920 3010
rect 24180 1810 25780 3010
<< ndiff >>
rect 32180 2780 33780 2810
rect 32180 1640 32210 2780
rect 33750 1640 33780 2780
rect 32180 1610 33780 1640
rect 35380 2780 36980 2810
rect 35380 1640 35410 2780
rect 36950 1640 36980 2780
rect 35380 1610 36980 1640
rect 37040 2780 38640 2810
rect 37040 1640 37070 2780
rect 38610 1640 38640 2780
rect 37040 1610 38640 1640
rect 40240 2780 41840 2810
rect 40240 1640 40270 2780
rect 41810 1640 41840 2780
rect 40240 1610 41840 1640
rect 43440 2780 45040 2810
rect 43440 1640 43470 2780
rect 45010 1640 45040 2780
rect 43440 1610 45040 1640
rect 46640 2780 48240 2810
rect 46640 1640 46670 2780
rect 48210 1640 48240 2780
rect 46640 1610 48240 1640
rect 49840 2780 51440 2810
rect 49840 1640 49870 2780
rect 51410 1640 51440 2780
rect 49840 1610 51440 1640
rect 51500 2780 53100 2810
rect 51500 1640 51530 2780
rect 53070 1640 53100 2780
rect 51500 1610 53100 1640
rect 54700 2780 56300 2810
rect 54700 1640 54730 2780
rect 56270 1640 56300 2780
rect 54700 1610 56300 1640
rect 57900 2780 59500 2810
rect 57900 1640 57930 2780
rect 59470 1640 59500 2780
rect 57900 1610 59500 1640
rect -4800 1170 -3200 1200
rect -4800 30 -4770 1170
rect -3230 30 -3200 1170
rect -4800 0 -3200 30
rect -1600 1170 0 1200
rect -1600 30 -1570 1170
rect -30 30 0 1170
rect -1600 0 0 30
rect 1600 1170 3200 1200
rect 1600 30 1630 1170
rect 3170 30 3200 1170
rect 1600 0 3200 30
rect 3260 1170 4860 1200
rect 3260 30 3290 1170
rect 4830 30 4860 1170
rect 3260 0 4860 30
rect 6460 1170 8060 1200
rect 6460 30 6490 1170
rect 8030 30 8060 1170
rect 6460 0 8060 30
rect 9660 1170 11260 1200
rect 9660 30 9690 1170
rect 11230 30 11260 1170
rect 9660 0 11260 30
rect 11320 1170 12920 1200
rect 11320 30 11350 1170
rect 12890 30 12920 1170
rect 11320 0 12920 30
rect 14520 1170 16120 1200
rect 14520 30 14550 1170
rect 16090 30 16120 1170
rect 14520 0 16120 30
rect 17720 1170 19320 1200
rect 17720 30 17750 1170
rect 19290 30 19320 1170
rect 17720 0 19320 30
rect 19380 1170 20980 1200
rect 19380 30 19410 1170
rect 20950 30 20980 1170
rect 19380 0 20980 30
rect 22580 1170 24180 1200
rect 22580 30 22610 1170
rect 24150 30 24180 1170
rect 22580 0 24180 30
rect 25780 1170 27380 1200
rect 25780 30 25810 1170
rect 27350 30 27380 1170
rect 25780 0 27380 30
rect 28980 1170 30580 1200
rect 28980 30 29010 1170
rect 30550 30 30580 1170
rect 28980 0 30580 30
rect 32180 1170 33780 1200
rect 32180 30 32210 1170
rect 33750 30 33780 1170
rect 32180 0 33780 30
rect 35380 1170 36980 1200
rect 35380 30 35410 1170
rect 36950 30 36980 1170
rect 35380 0 36980 30
rect 38580 1170 40180 1200
rect 38580 30 38610 1170
rect 40150 30 40180 1170
rect 38580 0 40180 30
rect 40240 1170 41840 1200
rect 40240 30 40270 1170
rect 41810 30 41840 1170
rect 40240 0 41840 30
rect 43440 1170 45040 1200
rect 43440 30 43470 1170
rect 45010 30 45040 1170
rect 43440 0 45040 30
rect 46640 1170 48240 1200
rect 46640 30 46670 1170
rect 48210 30 48240 1170
rect 46640 0 48240 30
rect 48300 1170 49900 1200
rect 48300 30 48330 1170
rect 49870 30 49900 1170
rect 48300 0 49900 30
rect 51500 1170 53100 1200
rect 51500 30 51530 1170
rect 53070 30 53100 1170
rect 51500 0 53100 30
rect 54700 1170 56300 1200
rect 54700 30 54730 1170
rect 56270 30 56300 1170
rect 54700 0 56300 30
rect 56360 1170 57960 1200
rect 56360 30 56390 1170
rect 57930 30 57960 1170
rect 56360 0 57960 30
rect 59560 1170 61160 1200
rect 59560 30 59590 1170
rect 61130 30 61160 1170
rect 59560 0 61160 30
rect 62760 1170 64360 1200
rect 62760 30 62790 1170
rect 64330 30 64360 1170
rect 62760 0 64360 30
<< pdiff >>
rect -3260 4520 -1660 4550
rect -3260 3380 -3230 4520
rect -1690 3380 -1660 4520
rect -3260 3350 -1660 3380
rect -60 4520 1540 4550
rect -60 3380 -30 4520
rect 1510 3380 1540 4520
rect -60 3350 1540 3380
rect 3140 4520 4740 4550
rect 3140 3380 3170 4520
rect 4710 3380 4740 4520
rect 3140 3350 4740 3380
rect 4800 4520 6400 4550
rect 4800 3380 4830 4520
rect 6370 3380 6400 4520
rect 4800 3350 6400 3380
rect 8000 4520 9600 4550
rect 8000 3380 8030 4520
rect 9570 3380 9600 4520
rect 8000 3350 9600 3380
rect 11200 4520 12800 4550
rect 11200 3380 11230 4520
rect 12770 3380 12800 4520
rect 11200 3350 12800 3380
rect 12860 4520 14460 4550
rect 12860 3380 12890 4520
rect 14430 3380 14460 4520
rect 12860 3350 14460 3380
rect 16060 4520 17660 4550
rect 16060 3380 16090 4520
rect 17630 3380 17660 4520
rect 16060 3350 17660 3380
rect 19260 4520 20860 4550
rect 19260 3380 19290 4520
rect 20830 3380 20860 4520
rect 19260 3350 20860 3380
rect 20920 4520 22520 4550
rect 20920 3380 20950 4520
rect 22490 3380 22520 4520
rect 20920 3350 22520 3380
rect 24120 4520 25720 4550
rect 24120 3380 24150 4520
rect 25690 3380 25720 4520
rect 24120 3350 25720 3380
rect 27320 4520 28920 4550
rect 27320 3380 27350 4520
rect 28890 3380 28920 4520
rect 27320 3350 28920 3380
rect 30520 4520 32120 4550
rect 30520 3380 30550 4520
rect 32090 3380 32120 4520
rect 30520 3350 32120 3380
rect 33720 4520 35320 4550
rect 33720 3380 33750 4520
rect 35290 3380 35320 4520
rect 33720 3350 35320 3380
rect 36920 4520 38520 4550
rect 36920 3380 36950 4520
rect 38490 3380 38520 4520
rect 36920 3350 38520 3380
rect 40120 4520 41720 4550
rect 40120 3380 40150 4520
rect 41690 3380 41720 4520
rect 40120 3350 41720 3380
rect 41780 4520 43380 4550
rect 41780 3380 41810 4520
rect 43350 3380 43380 4520
rect 41780 3350 43380 3380
rect 44980 4520 46580 4550
rect 44980 3380 45010 4520
rect 46550 3380 46580 4520
rect 44980 3350 46580 3380
rect 48180 4520 49780 4550
rect 48180 3380 48210 4520
rect 49750 3380 49780 4520
rect 48180 3350 49780 3380
rect 49840 4520 51440 4550
rect 49840 3380 49870 4520
rect 51410 3380 51440 4520
rect 49840 3350 51440 3380
rect 53040 4520 54640 4550
rect 53040 3380 53070 4520
rect 54610 3380 54640 4520
rect 53040 3350 54640 3380
rect 56240 4520 57840 4550
rect 56240 3380 56270 4520
rect 57810 3380 57840 4520
rect 56240 3350 57840 3380
rect 57900 4520 59500 4550
rect 57900 3380 57930 4520
rect 59470 3380 59500 4520
rect 57900 3350 59500 3380
rect 61100 4520 62700 4550
rect 61100 3380 61130 4520
rect 62670 3380 62700 4520
rect 61100 3350 62700 3380
rect 64300 4520 65900 4550
rect 64300 3380 64330 4520
rect 65870 3380 65900 4520
rect 64300 3350 65900 3380
rect -3260 2980 -1660 3010
rect -3260 1840 -3230 2980
rect -1690 1840 -1660 2980
rect -3260 1810 -1660 1840
rect -60 2980 1540 3010
rect -60 1840 -30 2980
rect 1510 1840 1540 2980
rect -60 1810 1540 1840
rect 3140 2980 4740 3010
rect 3140 1840 3170 2980
rect 4710 1840 4740 2980
rect 3140 1810 4740 1840
rect 4800 2980 6400 3010
rect 4800 1840 4830 2980
rect 6370 1840 6400 2980
rect 4800 1810 6400 1840
rect 8000 2980 9600 3010
rect 8000 1840 8030 2980
rect 9570 1840 9600 2980
rect 8000 1810 9600 1840
rect 9660 2980 11260 3010
rect 9660 1840 9690 2980
rect 11230 1840 11260 2980
rect 9660 1810 11260 1840
rect 12860 2980 14460 3010
rect 12860 1840 12890 2980
rect 14430 1840 14460 2980
rect 12860 1810 14460 1840
rect 16060 2980 17660 3010
rect 16060 1840 16090 2980
rect 17630 1840 17660 2980
rect 16060 1810 17660 1840
rect 17720 2980 19320 3010
rect 17720 1840 17750 2980
rect 19290 1840 19320 2980
rect 17720 1810 19320 1840
rect 20920 2980 22520 3010
rect 20920 1840 20950 2980
rect 22490 1840 22520 2980
rect 20920 1810 22520 1840
rect 22580 2980 24180 3010
rect 22580 1840 22610 2980
rect 24150 1840 24180 2980
rect 22580 1810 24180 1840
rect 25780 2980 27380 3010
rect 25780 1840 25810 2980
rect 27350 1840 27380 2980
rect 25780 1810 27380 1840
<< ndiffc >>
rect 32210 1640 33750 2780
rect 35410 1640 36950 2780
rect 37070 1640 38610 2780
rect 40270 1640 41810 2780
rect 43470 1640 45010 2780
rect 46670 1640 48210 2780
rect 49870 1640 51410 2780
rect 51530 1640 53070 2780
rect 54730 1640 56270 2780
rect 57930 1640 59470 2780
rect -4770 30 -3230 1170
rect -1570 30 -30 1170
rect 1630 30 3170 1170
rect 3290 30 4830 1170
rect 6490 30 8030 1170
rect 9690 30 11230 1170
rect 11350 30 12890 1170
rect 14550 30 16090 1170
rect 17750 30 19290 1170
rect 19410 30 20950 1170
rect 22610 30 24150 1170
rect 25810 30 27350 1170
rect 29010 30 30550 1170
rect 32210 30 33750 1170
rect 35410 30 36950 1170
rect 38610 30 40150 1170
rect 40270 30 41810 1170
rect 43470 30 45010 1170
rect 46670 30 48210 1170
rect 48330 30 49870 1170
rect 51530 30 53070 1170
rect 54730 30 56270 1170
rect 56390 30 57930 1170
rect 59590 30 61130 1170
rect 62790 30 64330 1170
<< pdiffc >>
rect -3230 3380 -1690 4520
rect -30 3380 1510 4520
rect 3170 3380 4710 4520
rect 4830 3380 6370 4520
rect 8030 3380 9570 4520
rect 11230 3380 12770 4520
rect 12890 3380 14430 4520
rect 16090 3380 17630 4520
rect 19290 3380 20830 4520
rect 20950 3380 22490 4520
rect 24150 3380 25690 4520
rect 27350 3380 28890 4520
rect 30550 3380 32090 4520
rect 33750 3380 35290 4520
rect 36950 3380 38490 4520
rect 40150 3380 41690 4520
rect 41810 3380 43350 4520
rect 45010 3380 46550 4520
rect 48210 3380 49750 4520
rect 49870 3380 51410 4520
rect 53070 3380 54610 4520
rect 56270 3380 57810 4520
rect 57930 3380 59470 4520
rect 61130 3380 62670 4520
rect 64330 3380 65870 4520
rect -3230 1840 -1690 2980
rect -30 1840 1510 2980
rect 3170 1840 4710 2980
rect 4830 1840 6370 2980
rect 8030 1840 9570 2980
rect 9690 1840 11230 2980
rect 12890 1840 14430 2980
rect 16090 1840 17630 2980
rect 17750 1840 19290 2980
rect 20950 1840 22490 2980
rect 22610 1840 24150 2980
rect 25810 1840 27350 2980
<< psubdiff >>
rect 59500 2780 61100 2810
rect 59500 1640 59530 2780
rect 61070 1640 61100 2780
rect 59500 1610 61100 1640
rect -6400 1170 -4800 1200
rect -6400 30 -6370 1170
rect -4830 30 -4800 1170
rect -6400 0 -4800 30
rect 64360 1170 65960 1200
rect 64360 30 64390 1170
rect 65930 30 65960 1170
rect 64360 0 65960 30
<< nsubdiff >>
rect -4860 4520 -3260 4550
rect -4860 3380 -4830 4520
rect -3290 3380 -3260 4520
rect -4860 3350 -3260 3380
rect 65900 4520 67500 4550
rect 65900 3380 65930 4520
rect 67470 3380 67500 4520
rect 65900 3350 67500 3380
rect -4860 2980 -3260 3010
rect -4860 1840 -4830 2980
rect -3290 1840 -3260 2980
rect -4860 1810 -3260 1840
<< psubdiffcont >>
rect 59530 1640 61070 2780
rect -6370 30 -4830 1170
rect 64390 30 65930 1170
<< nsubdiffcont >>
rect -4830 3380 -3290 4520
rect 65930 3380 67470 4520
rect -4830 1840 -3290 2980
<< poly >>
rect 14910 4930 15000 4950
rect 14910 4890 14930 4930
rect 14980 4890 15000 4930
rect 14910 4880 15000 4890
rect 23090 4930 23180 4950
rect 23090 4890 23110 4930
rect 23160 4890 23180 4930
rect 23090 4880 23180 4890
rect 39460 4930 39550 4940
rect 39460 4890 39480 4930
rect 39530 4890 39550 4930
rect 39460 4880 39550 4890
rect 47640 4930 47730 4940
rect 47640 4890 47660 4930
rect 47710 4890 47730 4930
rect 47640 4880 47730 4890
rect -1620 4680 -1530 4700
rect -1620 4640 -1600 4680
rect -1550 4640 -1530 4680
rect -1620 4630 -1530 4640
rect 1580 4680 1670 4700
rect 1580 4640 1600 4680
rect 1650 4640 1670 4680
rect 1580 4630 1670 4640
rect 6440 4680 6530 4700
rect 6440 4640 6460 4680
rect 6510 4640 6530 4680
rect 6440 4630 6530 4640
rect 9640 4680 9730 4700
rect 9640 4640 9660 4680
rect 9710 4640 9730 4680
rect 9640 4630 9730 4640
rect 13210 4680 13300 4700
rect 13210 4640 13230 4680
rect 13280 4660 13300 4680
rect 13510 4680 13600 4700
rect 13510 4660 13530 4680
rect 13280 4640 13530 4660
rect 13580 4640 13600 4680
rect 13210 4630 13600 4640
rect -1610 4580 -1580 4630
rect 1590 4580 1620 4630
rect 6450 4580 6480 4630
rect 9650 4580 9680 4630
rect 14940 4580 14970 4880
rect 17700 4680 17790 4700
rect 17700 4640 17720 4680
rect 17770 4640 17790 4680
rect 17700 4630 17790 4640
rect 21150 4680 21240 4700
rect 21150 4640 21170 4680
rect 21220 4660 21240 4680
rect 21450 4680 21540 4700
rect 21450 4660 21470 4680
rect 21220 4640 21470 4660
rect 21520 4640 21540 4680
rect 21150 4630 21540 4640
rect 17710 4580 17740 4630
rect 23120 4580 23150 4880
rect 25760 4680 25850 4700
rect 25760 4640 25780 4680
rect 25830 4640 25850 4680
rect 25760 4630 25850 4640
rect 28960 4680 29050 4700
rect 28960 4640 28980 4680
rect 29030 4640 29050 4680
rect 28960 4630 29050 4640
rect 33590 4680 33680 4700
rect 33590 4640 33610 4680
rect 33660 4640 33680 4680
rect 33590 4630 33680 4640
rect 36790 4680 36880 4700
rect 36790 4640 36810 4680
rect 36860 4640 36880 4680
rect 36790 4630 36880 4640
rect 25770 4580 25810 4630
rect 28970 4580 29010 4630
rect 33630 4580 33670 4630
rect 36830 4580 36870 4630
rect 39490 4580 39520 4880
rect 41100 4680 41190 4700
rect 41100 4640 41120 4680
rect 41170 4660 41190 4680
rect 41400 4680 41490 4700
rect 41400 4660 41420 4680
rect 41170 4640 41420 4660
rect 41470 4640 41490 4680
rect 41100 4630 41490 4640
rect 44850 4680 44940 4700
rect 44850 4640 44870 4680
rect 44920 4640 44940 4680
rect 44850 4630 44940 4640
rect 44900 4580 44930 4630
rect 47670 4580 47700 4880
rect 67430 4800 67520 4820
rect 67430 4760 67450 4800
rect 67500 4780 67520 4800
rect 67770 4800 67860 4820
rect 67770 4780 67790 4800
rect 67500 4760 67790 4780
rect 67840 4760 67860 4800
rect 67430 4750 67860 4760
rect 49040 4680 49130 4700
rect 49040 4640 49060 4680
rect 49110 4660 49130 4680
rect 49340 4680 49430 4700
rect 49340 4660 49360 4680
rect 49110 4640 49360 4660
rect 49410 4640 49430 4680
rect 49040 4630 49430 4640
rect 52910 4680 53000 4700
rect 52910 4640 52930 4680
rect 52980 4640 53000 4680
rect 52910 4630 53000 4640
rect 56110 4680 56200 4700
rect 56110 4640 56130 4680
rect 56180 4640 56200 4680
rect 56110 4630 56200 4640
rect 60970 4680 61060 4700
rect 60970 4640 60990 4680
rect 61040 4640 61060 4680
rect 60970 4630 61060 4640
rect 64170 4680 64260 4700
rect 64170 4640 64190 4680
rect 64240 4640 64260 4680
rect 64170 4630 64260 4640
rect 52960 4580 52990 4630
rect 56160 4580 56190 4630
rect 61020 4580 61050 4630
rect 64220 4580 64250 4630
rect -1660 4550 -60 4580
rect 1540 4550 3140 4580
rect 6400 4550 8000 4580
rect 9600 4550 11200 4580
rect 14460 4550 16060 4580
rect 17660 4550 19260 4580
rect 22520 4550 24120 4580
rect 25720 4550 27320 4580
rect 28920 4550 30520 4580
rect 32120 4550 33720 4580
rect 35320 4550 36920 4580
rect 38520 4550 40120 4580
rect 43380 4550 44980 4580
rect 46580 4550 48180 4580
rect 51440 4550 53040 4580
rect 54640 4550 56240 4580
rect 59500 4550 61100 4580
rect 62700 4550 64300 4580
rect -1660 3320 -60 3350
rect 1540 3320 3140 3350
rect 6400 3320 8000 3350
rect 9600 3320 11200 3350
rect 14460 3320 16060 3350
rect 17660 3320 19260 3350
rect 22520 3320 24120 3350
rect 25720 3320 27320 3350
rect 28920 3320 30520 3350
rect 32120 3320 33720 3350
rect 35320 3320 36920 3350
rect 38520 3320 40120 3350
rect 43380 3320 44980 3350
rect 46580 3320 48180 3350
rect 51440 3320 53040 3350
rect 54640 3320 56240 3350
rect 59500 3320 61100 3350
rect 62700 3320 64300 3350
rect -1610 3140 -1520 3160
rect -1610 3100 -1590 3140
rect -1540 3100 -1520 3140
rect -1610 3090 -1520 3100
rect 3050 3140 3140 3160
rect 3050 3100 3070 3140
rect 3120 3100 3140 3140
rect 3050 3090 3140 3100
rect 5700 3140 5790 3160
rect 5700 3100 5720 3140
rect 5770 3120 5790 3140
rect 6000 3140 6090 3160
rect 6000 3120 6020 3140
rect 5770 3100 6020 3120
rect 6070 3100 6090 3140
rect 5700 3090 6090 3100
rect 7910 3140 8000 3160
rect 7910 3100 7930 3140
rect 7980 3100 8000 3140
rect 7910 3090 8000 3100
rect 9910 3140 10000 3160
rect 9910 3100 9930 3140
rect 9980 3120 10000 3140
rect 10210 3140 10300 3160
rect 10210 3120 10230 3140
rect 9980 3100 10230 3120
rect 10280 3100 10300 3140
rect 9910 3090 10300 3100
rect 12770 3140 12860 3160
rect 12770 3100 12790 3140
rect 12840 3100 12860 3140
rect 12770 3090 12860 3100
rect -1600 3040 -1570 3090
rect 3110 3040 3140 3090
rect 7970 3040 8000 3090
rect 12830 3040 12860 3090
rect -1660 3010 -60 3040
rect 1540 3010 3140 3040
rect 6400 3010 8000 3040
rect 11260 3010 12860 3040
rect 14460 3140 14550 3160
rect 14460 3100 14480 3140
rect 14530 3100 14550 3140
rect 14460 3090 14550 3100
rect 17020 3140 17110 3160
rect 17020 3100 17040 3140
rect 17090 3120 17110 3140
rect 17320 3140 17410 3160
rect 17320 3120 17340 3140
rect 17090 3100 17340 3120
rect 17390 3100 17410 3140
rect 17020 3090 17410 3100
rect 19320 3140 19410 3160
rect 19320 3100 19340 3140
rect 19390 3100 19410 3140
rect 19320 3090 19410 3100
rect 21230 3140 21320 3160
rect 21230 3100 21250 3140
rect 21300 3120 21320 3140
rect 21530 3140 21620 3160
rect 21530 3120 21550 3140
rect 21300 3100 21550 3120
rect 21600 3100 21620 3140
rect 21230 3090 21620 3100
rect 24180 3140 24270 3160
rect 24180 3100 24200 3140
rect 24250 3100 24270 3140
rect 24180 3090 24270 3100
rect 14460 3040 14490 3090
rect 19320 3040 19350 3090
rect 24180 3040 24210 3090
rect 14460 3010 16060 3040
rect 19320 3010 20920 3040
rect 24180 3010 25780 3040
rect 43250 2970 43750 2990
rect 43250 2930 43270 2970
rect 43320 2960 43680 2970
rect 43320 2930 43340 2960
rect 43250 2920 43340 2930
rect 43660 2930 43680 2960
rect 43730 2930 43750 2970
rect 43660 2920 43750 2930
rect 33780 2810 35380 2840
rect 38640 2810 40240 2840
rect 41840 2810 43440 2840
rect 45040 2810 46640 2840
rect 48240 2810 49840 2840
rect 53100 2810 54700 2840
rect 56300 2810 57900 2840
rect -1660 1780 -60 1810
rect 1540 1780 3140 1810
rect 6400 1780 8000 1810
rect 11260 1780 12860 1810
rect 14460 1780 16060 1810
rect 19320 1780 20920 1810
rect 24180 1780 25780 1810
rect 13490 1690 13580 1710
rect 13490 1650 13510 1690
rect 13560 1670 13580 1690
rect 13860 1690 13950 1710
rect 13860 1670 13880 1690
rect 13560 1650 13880 1670
rect 13930 1650 13950 1690
rect 13490 1640 13950 1650
rect 33780 1580 35380 1610
rect 38640 1580 40240 1610
rect 41840 1580 43440 1610
rect 45040 1580 46640 1610
rect 48240 1580 49840 1610
rect 53100 1580 54700 1610
rect 56300 1580 57900 1610
rect 13490 1560 13580 1580
rect 13490 1520 13510 1560
rect 13560 1540 13580 1560
rect 13860 1560 13950 1580
rect 13860 1540 13880 1560
rect 13560 1520 13880 1540
rect 13930 1520 13950 1560
rect 13490 1510 13950 1520
rect 18100 1560 18190 1580
rect 18100 1520 18120 1560
rect 18170 1540 18190 1560
rect 18430 1560 18520 1580
rect 18430 1540 18450 1560
rect 18170 1520 18450 1540
rect 18500 1520 18520 1560
rect 18100 1510 18520 1520
rect 33780 1570 33870 1580
rect 33780 1530 33800 1570
rect 33850 1530 33870 1570
rect 33780 1510 33870 1530
rect 38640 1570 38730 1580
rect 38640 1530 38660 1570
rect 38710 1530 38730 1570
rect 38640 1510 38730 1530
rect 41840 1570 41930 1580
rect 41840 1530 41860 1570
rect 41910 1530 41930 1570
rect 41840 1510 41930 1530
rect 46550 1570 46640 1580
rect 46550 1530 46570 1570
rect 46620 1530 46640 1570
rect 46550 1510 46640 1530
rect 49750 1570 49840 1580
rect 49750 1530 49770 1570
rect 49820 1530 49840 1570
rect 49750 1510 49840 1530
rect 54610 1570 54700 1580
rect 54610 1530 54630 1570
rect 54680 1530 54700 1570
rect 54610 1510 54700 1530
rect 57760 1570 57850 1580
rect 57760 1530 57780 1570
rect 57830 1530 57850 1570
rect 57760 1510 57850 1530
rect 12920 1440 13010 1460
rect 12920 1400 12940 1440
rect 12990 1400 13010 1440
rect 12920 1390 13010 1400
rect 13490 1440 13580 1460
rect 13490 1400 13510 1440
rect 13560 1420 13580 1440
rect 13860 1440 13950 1460
rect 13860 1420 13880 1440
rect 13560 1400 13880 1420
rect 13930 1400 13950 1440
rect 13490 1390 13950 1400
rect 20980 1440 21070 1460
rect 20980 1400 21000 1440
rect 21050 1400 21070 1440
rect 20980 1390 21070 1400
rect 38490 1440 38580 1460
rect 38490 1400 38510 1440
rect 38560 1400 38580 1440
rect 38490 1390 38580 1400
rect 46550 1440 46640 1460
rect 46550 1400 46570 1440
rect 46620 1400 46640 1440
rect 46550 1390 46640 1400
rect 0 1330 90 1350
rect 0 1290 20 1330
rect 70 1290 90 1330
rect 0 1280 90 1290
rect 4860 1330 4950 1350
rect 4860 1290 4880 1330
rect 4930 1290 4950 1330
rect 4860 1280 4950 1290
rect 8060 1330 8150 1350
rect 8060 1290 8080 1330
rect 8130 1290 8150 1330
rect 8060 1280 8150 1290
rect 11180 1330 11270 1350
rect 11180 1290 11200 1330
rect 11250 1310 11270 1330
rect 11480 1330 11570 1350
rect 11480 1310 11500 1330
rect 11250 1290 11500 1310
rect 11550 1290 11570 1330
rect 11180 1280 11570 1290
rect 0 1230 30 1280
rect 4860 1230 4890 1280
rect 8060 1230 8090 1280
rect 12920 1230 12950 1390
rect 16120 1330 16210 1350
rect 16120 1290 16140 1330
rect 16190 1290 16210 1330
rect 16120 1280 16210 1290
rect 19240 1330 19330 1350
rect 19240 1290 19260 1330
rect 19310 1310 19330 1330
rect 19540 1330 19630 1350
rect 19540 1310 19560 1330
rect 19310 1290 19560 1310
rect 19610 1290 19630 1330
rect 19240 1280 19630 1290
rect 16120 1230 16150 1280
rect 20980 1230 21010 1390
rect 24180 1330 24270 1350
rect 24180 1290 24200 1330
rect 24250 1290 24270 1330
rect 24180 1280 24270 1290
rect 27380 1330 27470 1350
rect 27380 1290 27400 1330
rect 27450 1290 27470 1330
rect 27380 1280 27470 1290
rect 32090 1330 32180 1350
rect 32090 1290 32110 1330
rect 32160 1290 32180 1330
rect 32090 1280 32180 1290
rect 35290 1330 35380 1350
rect 35290 1290 35310 1330
rect 35360 1290 35380 1330
rect 35290 1280 35380 1290
rect 24180 1230 24210 1280
rect 27380 1230 27410 1280
rect 32150 1230 32180 1280
rect 35350 1230 35380 1280
rect 38550 1230 38580 1390
rect 39930 1330 40020 1350
rect 39930 1290 39950 1330
rect 40000 1310 40020 1330
rect 40230 1330 40320 1350
rect 40230 1310 40250 1330
rect 40000 1290 40250 1310
rect 40300 1290 40320 1330
rect 39930 1280 40320 1290
rect 43350 1330 43440 1350
rect 43350 1290 43370 1330
rect 43420 1290 43440 1330
rect 43350 1280 43440 1290
rect 43410 1230 43440 1280
rect 46610 1230 46640 1390
rect 47990 1330 48080 1350
rect 47990 1290 48010 1330
rect 48060 1310 48080 1330
rect 48290 1330 48380 1350
rect 48290 1310 48310 1330
rect 48060 1290 48310 1310
rect 48360 1290 48380 1330
rect 47990 1280 48380 1290
rect 51410 1330 51500 1350
rect 51410 1290 51430 1330
rect 51480 1290 51500 1330
rect 51410 1280 51500 1290
rect 54610 1330 54700 1350
rect 54610 1290 54630 1330
rect 54680 1290 54700 1330
rect 54610 1280 54700 1290
rect 59470 1330 59560 1350
rect 59470 1290 59490 1330
rect 59540 1290 59560 1330
rect 59470 1280 59560 1290
rect 51470 1230 51500 1280
rect 54670 1230 54700 1280
rect 59530 1230 59560 1280
rect -3200 1200 -1600 1230
rect 0 1200 1600 1230
rect 4860 1200 6460 1230
rect 8060 1200 9660 1230
rect 12920 1200 14520 1230
rect 16120 1200 17720 1230
rect 20980 1200 22580 1230
rect 24180 1200 25780 1230
rect 27380 1200 28980 1230
rect 30580 1200 32180 1230
rect 33780 1200 35380 1230
rect 36980 1200 38580 1230
rect 41840 1200 43440 1230
rect 45040 1200 46640 1230
rect 49900 1200 51500 1230
rect 53100 1200 54700 1230
rect 57960 1200 59560 1230
rect 61160 1200 62760 1230
rect -3200 -30 -1600 0
rect 0 -30 1600 0
rect 4860 -30 6460 0
rect 8060 -30 9660 0
rect 12920 -30 14520 0
rect 16120 -30 17720 0
rect 20980 -30 22580 0
rect 24180 -30 25780 0
rect 27380 -30 28980 0
rect 30580 -30 32180 0
rect 33780 -30 35380 0
rect 36980 -30 38580 0
rect 41840 -30 43440 0
rect 45040 -30 46640 0
rect 49900 -30 51500 0
rect 53100 -30 54700 0
rect 57960 -30 59560 0
rect 61160 -30 62760 0
rect -3200 -40 -3110 -30
rect -3200 -80 -3180 -40
rect -3130 -80 -3110 -40
rect -3200 -100 -3110 -80
rect 62670 -40 62760 -30
rect 62670 -80 62690 -40
rect 62740 -80 62760 -40
rect 62670 -100 62760 -80
<< polycont >>
rect 14930 4890 14980 4930
rect 23110 4890 23160 4930
rect 39480 4890 39530 4930
rect 47660 4890 47710 4930
rect -1600 4640 -1550 4680
rect 1600 4640 1650 4680
rect 6460 4640 6510 4680
rect 9660 4640 9710 4680
rect 13230 4640 13280 4680
rect 13530 4640 13580 4680
rect 17720 4640 17770 4680
rect 21170 4640 21220 4680
rect 21470 4640 21520 4680
rect 25780 4640 25830 4680
rect 28980 4640 29030 4680
rect 33610 4640 33660 4680
rect 36810 4640 36860 4680
rect 41120 4640 41170 4680
rect 41420 4640 41470 4680
rect 44870 4640 44920 4680
rect 67450 4760 67500 4800
rect 67790 4760 67840 4800
rect 49060 4640 49110 4680
rect 49360 4640 49410 4680
rect 52930 4640 52980 4680
rect 56130 4640 56180 4680
rect 60990 4640 61040 4680
rect 64190 4640 64240 4680
rect -1590 3100 -1540 3140
rect 3070 3100 3120 3140
rect 5720 3100 5770 3140
rect 6020 3100 6070 3140
rect 7930 3100 7980 3140
rect 9930 3100 9980 3140
rect 10230 3100 10280 3140
rect 12790 3100 12840 3140
rect 14480 3100 14530 3140
rect 17040 3100 17090 3140
rect 17340 3100 17390 3140
rect 19340 3100 19390 3140
rect 21250 3100 21300 3140
rect 21550 3100 21600 3140
rect 24200 3100 24250 3140
rect 43270 2930 43320 2970
rect 43680 2930 43730 2970
rect 13510 1650 13560 1690
rect 13880 1650 13930 1690
rect 13510 1520 13560 1560
rect 13880 1520 13930 1560
rect 18120 1520 18170 1560
rect 18450 1520 18500 1560
rect 33800 1530 33850 1570
rect 38660 1530 38710 1570
rect 41860 1530 41910 1570
rect 46570 1530 46620 1570
rect 49770 1530 49820 1570
rect 54630 1530 54680 1570
rect 57780 1530 57830 1570
rect 12940 1400 12990 1440
rect 13510 1400 13560 1440
rect 13880 1400 13930 1440
rect 21000 1400 21050 1440
rect 38510 1400 38560 1440
rect 46570 1400 46620 1440
rect 20 1290 70 1330
rect 4880 1290 4930 1330
rect 8080 1290 8130 1330
rect 11200 1290 11250 1330
rect 11500 1290 11550 1330
rect 16140 1290 16190 1330
rect 19260 1290 19310 1330
rect 19560 1290 19610 1330
rect 24200 1290 24250 1330
rect 27400 1290 27450 1330
rect 32110 1290 32160 1330
rect 35310 1290 35360 1330
rect 39950 1290 40000 1330
rect 40250 1290 40300 1330
rect 43370 1290 43420 1330
rect 48010 1290 48060 1330
rect 48310 1290 48360 1330
rect 51430 1290 51480 1330
rect 54630 1290 54680 1330
rect 59490 1290 59540 1330
rect -3180 -80 -3130 -40
rect 62690 -80 62740 -40
<< locali >>
rect 14910 4930 15000 4950
rect 14910 4920 14930 4930
rect 13380 4890 14930 4920
rect 14980 4920 15000 4930
rect 23090 4930 23180 4950
rect 23090 4920 23110 4930
rect 14980 4890 23110 4920
rect 23160 4920 23180 4930
rect 39460 4930 39550 4940
rect 39460 4920 39480 4930
rect 23160 4890 39480 4920
rect 39530 4920 39550 4930
rect 47640 4930 47730 4940
rect 47640 4920 47660 4930
rect 39530 4890 47660 4920
rect 47710 4920 47730 4930
rect 47710 4890 67890 4920
rect 13380 4880 67890 4890
rect -1620 4680 -1530 4700
rect -1620 4670 -1600 4680
rect -1710 4640 -1600 4670
rect -1550 4640 -1530 4680
rect -1710 4630 -1530 4640
rect 1580 4680 1670 4700
rect 1580 4640 1600 4680
rect 1650 4670 1670 4680
rect 6440 4680 6530 4700
rect 6440 4670 6460 4680
rect 1650 4640 6460 4670
rect 6510 4670 6530 4680
rect 9640 4680 9730 4700
rect 9640 4670 9660 4680
rect 6510 4640 9660 4670
rect 9710 4670 9730 4680
rect 13210 4680 13300 4700
rect 13210 4670 13230 4680
rect 9710 4640 13230 4670
rect 13280 4640 13300 4680
rect 1580 4630 13300 4640
rect -1710 4540 -1670 4630
rect 11210 4540 11250 4630
rect 13380 4540 13420 4880
rect 13510 4680 13600 4700
rect 13510 4640 13530 4680
rect 13580 4670 13600 4680
rect 17700 4680 17790 4700
rect 17700 4670 17720 4680
rect 13580 4640 17720 4670
rect 17770 4670 17790 4680
rect 21150 4680 21240 4700
rect 21150 4670 21170 4680
rect 17770 4640 21170 4670
rect 21220 4640 21240 4680
rect 13510 4630 21240 4640
rect 19270 4540 19310 4630
rect 21320 4540 21360 4880
rect 21450 4680 21540 4700
rect 21450 4640 21470 4680
rect 21520 4670 21540 4680
rect 25760 4680 25850 4700
rect 25760 4670 25780 4680
rect 21520 4640 25780 4670
rect 25830 4670 25850 4680
rect 28960 4680 29050 4700
rect 28960 4670 28980 4680
rect 25830 4640 28980 4670
rect 29030 4670 29050 4680
rect 33590 4680 33680 4700
rect 33590 4670 33610 4680
rect 29030 4640 33610 4670
rect 33660 4670 33680 4680
rect 36790 4680 36880 4700
rect 36790 4670 36810 4680
rect 33660 4640 36810 4670
rect 36860 4670 36880 4680
rect 41100 4680 41190 4700
rect 41100 4670 41120 4680
rect 36860 4640 41120 4670
rect 41170 4640 41190 4680
rect 21450 4630 41190 4640
rect 27330 4540 27370 4630
rect 35270 4540 35310 4630
rect 41280 4540 41320 4880
rect 41400 4680 41490 4700
rect 41400 4640 41420 4680
rect 41470 4670 41490 4680
rect 44850 4680 44940 4700
rect 44850 4670 44870 4680
rect 41470 4640 44870 4670
rect 44920 4670 44940 4680
rect 49040 4680 49130 4700
rect 49040 4670 49060 4680
rect 44920 4640 49060 4670
rect 49110 4640 49130 4680
rect 41400 4630 49130 4640
rect 43330 4540 43370 4630
rect 49220 4540 49260 4880
rect 67430 4800 67520 4820
rect 67430 4790 67450 4800
rect 61020 4760 67450 4790
rect 67500 4760 67520 4800
rect 61020 4750 67520 4760
rect 61020 4700 61060 4750
rect 49340 4680 49430 4700
rect 49340 4640 49360 4680
rect 49410 4670 49430 4680
rect 52910 4680 53000 4700
rect 52910 4670 52930 4680
rect 49410 4640 52930 4670
rect 52980 4670 53000 4680
rect 56110 4680 56200 4700
rect 56110 4670 56130 4680
rect 52980 4640 56130 4670
rect 56180 4670 56200 4680
rect 60970 4680 61060 4700
rect 60970 4670 60990 4680
rect 56180 4640 60990 4670
rect 61040 4640 61060 4680
rect 49340 4630 61060 4640
rect 64170 4680 64260 4700
rect 64170 4640 64190 4680
rect 64240 4670 64260 4680
rect 67480 4670 67520 4750
rect 64240 4640 64350 4670
rect 64170 4630 64350 4640
rect 67480 4630 67630 4670
rect 51390 4540 51430 4630
rect 64310 4540 64350 4630
rect -4850 4520 -1670 4540
rect -4850 3380 -4830 4520
rect -3290 3380 -3230 4520
rect -1690 3380 -1670 4520
rect -4850 3360 -1670 3380
rect -50 4520 1530 4540
rect -50 3380 -30 4520
rect 1510 3380 1530 4520
rect -50 3360 1530 3380
rect 3150 4520 4730 4540
rect 3150 3380 3170 4520
rect 4710 3380 4730 4520
rect 3150 3360 4730 3380
rect 4810 4520 6390 4540
rect 4810 3380 4830 4520
rect 6370 3380 6390 4520
rect 4810 3360 6390 3380
rect 8010 4520 9590 4540
rect 8010 3380 8030 4520
rect 9570 3380 9590 4520
rect 8010 3360 9590 3380
rect 11210 4520 12790 4540
rect 11210 3380 11230 4520
rect 12770 3380 12790 4520
rect 11210 3360 12790 3380
rect 12870 4520 14450 4540
rect 12870 3380 12890 4520
rect 14430 3380 14450 4520
rect 12870 3360 14450 3380
rect 16070 4520 17650 4540
rect 16070 3380 16090 4520
rect 17630 3380 17650 4520
rect 16070 3360 17650 3380
rect 19270 4520 20850 4540
rect 19270 3380 19290 4520
rect 20830 3380 20850 4520
rect 19270 3360 20850 3380
rect 20930 4520 22510 4540
rect 20930 3380 20950 4520
rect 22490 3380 22510 4520
rect 20930 3360 22510 3380
rect 24130 4520 25710 4540
rect 24130 3380 24150 4520
rect 25690 3380 25710 4520
rect 24130 3360 25710 3380
rect 27330 4520 28910 4540
rect 27330 3380 27350 4520
rect 28890 3380 28910 4520
rect 27330 3360 28910 3380
rect 30530 4520 32110 4540
rect 30530 3380 30550 4520
rect 32090 3380 32110 4520
rect 30530 3360 32110 3380
rect 33730 4520 35310 4540
rect 33730 3380 33750 4520
rect 35290 3380 35310 4520
rect 33730 3360 35310 3380
rect 36930 4520 38510 4540
rect 36930 3380 36950 4520
rect 38490 3380 38510 4520
rect 36930 3360 38510 3380
rect 40130 4520 41710 4540
rect 40130 3380 40150 4520
rect 41690 3380 41710 4520
rect 40130 3360 41710 3380
rect 41790 4520 43370 4540
rect 41790 3380 41810 4520
rect 43350 3380 43370 4520
rect 41790 3360 43370 3380
rect 44990 4520 46570 4540
rect 44990 3380 45010 4520
rect 46550 3380 46570 4520
rect 44990 3360 46570 3380
rect 48190 4520 49770 4540
rect 48190 3380 48210 4520
rect 49750 3380 49770 4520
rect 48190 3360 49770 3380
rect 49850 4520 51430 4540
rect 49850 3380 49870 4520
rect 51410 3380 51430 4520
rect 49850 3360 51430 3380
rect 53050 4520 54630 4540
rect 53050 3380 53070 4520
rect 54610 3380 54630 4520
rect 53050 3360 54630 3380
rect 56250 4520 57830 4540
rect 56250 3380 56270 4520
rect 57810 3380 57830 4520
rect 56250 3360 57830 3380
rect 57910 4520 59490 4540
rect 57910 3380 57930 4520
rect 59470 3380 59490 4520
rect 57910 3360 59490 3380
rect 61110 4520 62690 4540
rect 61110 3380 61130 4520
rect 62670 3380 62690 4520
rect 61110 3360 62690 3380
rect 64310 4520 67490 4540
rect 64310 3380 64330 4520
rect 65870 3380 65930 4520
rect 67470 3380 67490 4520
rect 64310 3360 67490 3380
rect 4690 3320 4730 3360
rect 9550 3320 9590 3360
rect 17610 3320 17650 3360
rect 24760 3320 24800 3360
rect 31340 3320 31380 3360
rect 37840 3320 37880 3360
rect 44990 3320 45030 3360
rect 53050 3320 53090 3360
rect 57910 3320 57950 3360
rect 4690 3280 57950 3320
rect -6460 3210 -1370 3250
rect -1410 3160 -1370 3210
rect -1610 3140 -1520 3160
rect -1610 3100 -1590 3140
rect -1540 3100 -1520 3140
rect -1410 3140 3140 3160
rect -1410 3120 3070 3140
rect -1610 3090 -1520 3100
rect 3050 3100 3070 3120
rect 3120 3130 3140 3140
rect 5700 3140 5790 3160
rect 5700 3130 5720 3140
rect 3120 3100 5720 3130
rect 5770 3100 5790 3140
rect 6000 3140 6090 3160
rect 3050 3090 5790 3100
rect -1710 3050 -1570 3090
rect -1710 3000 -1670 3050
rect 1490 3000 1530 3010
rect 5880 3000 5920 3120
rect 6000 3100 6020 3140
rect 6070 3130 6090 3140
rect 7910 3140 8000 3160
rect 7910 3130 7930 3140
rect 6070 3100 7930 3130
rect 7980 3130 8000 3140
rect 9910 3140 10000 3160
rect 9910 3130 9930 3140
rect 7980 3100 9930 3130
rect 9980 3100 10000 3140
rect 10210 3140 10300 3160
rect 6000 3090 10000 3100
rect 10100 3000 10140 3120
rect 10210 3100 10230 3140
rect 10280 3130 10300 3140
rect 12770 3140 12860 3160
rect 12770 3130 12790 3140
rect 10280 3100 12790 3130
rect 12840 3130 12860 3140
rect 14460 3140 14550 3160
rect 14460 3130 14480 3140
rect 12840 3100 14480 3130
rect 14530 3130 14550 3140
rect 17020 3140 17110 3160
rect 17020 3130 17040 3140
rect 14530 3100 17040 3130
rect 17090 3100 17110 3140
rect 17320 3140 17410 3160
rect 10210 3090 17110 3100
rect 17180 3000 17220 3120
rect 17320 3100 17340 3140
rect 17390 3130 17410 3140
rect 19320 3140 19410 3160
rect 19320 3130 19340 3140
rect 17390 3100 19340 3130
rect 19390 3130 19410 3140
rect 21230 3140 21320 3160
rect 21230 3130 21250 3140
rect 19390 3100 21250 3130
rect 21300 3100 21320 3140
rect 21530 3140 21620 3160
rect 17320 3090 21320 3100
rect 21400 3000 21440 3120
rect 21530 3100 21550 3140
rect 21600 3130 21620 3140
rect 24180 3140 24270 3160
rect 24180 3130 24200 3140
rect 21600 3100 24200 3130
rect 24250 3100 24270 3140
rect 21530 3090 24270 3100
rect 67590 3090 67630 4630
rect 43450 3050 67630 3090
rect 25790 3000 25830 3020
rect -4850 2980 -1670 3000
rect -4850 1840 -4830 2980
rect -3290 1840 -3230 2980
rect -1690 1840 -1670 2980
rect -4850 1820 -1670 1840
rect -50 2980 1530 3000
rect -50 1840 -30 2980
rect 1510 1840 1530 2980
rect -50 1820 1530 1840
rect 3150 2980 4730 3000
rect 3150 1840 3170 2980
rect 4710 1840 4730 2980
rect 3150 1820 4730 1840
rect 4810 2980 6390 3000
rect 4810 1840 4830 2980
rect 6370 1840 6390 2980
rect 4810 1820 6390 1840
rect 8010 2980 9590 3000
rect 8010 1840 8030 2980
rect 9570 1840 9590 2980
rect 8010 1820 9590 1840
rect 9670 2980 11250 3000
rect 9670 1840 9690 2980
rect 11230 1840 11250 2980
rect 9670 1820 11250 1840
rect 12870 2980 14450 3000
rect 12870 1840 12890 2980
rect 14430 1840 14450 2980
rect 12870 1820 14450 1840
rect 16070 2980 17650 3000
rect 16070 1840 16090 2980
rect 17630 1840 17650 2980
rect 16070 1820 17650 1840
rect 17730 2980 19310 3000
rect 17730 1840 17750 2980
rect 19290 1840 19310 2980
rect 17730 1820 19310 1840
rect 20930 2980 22510 3000
rect 20930 1840 20950 2980
rect 22490 1840 22510 2980
rect 20930 1820 22510 1840
rect 22590 2980 24170 3000
rect 22590 1840 22610 2980
rect 24150 1840 24170 2980
rect 22590 1820 24170 1840
rect 25790 2980 27370 3000
rect 25790 1840 25810 2980
rect 27350 1840 27370 2980
rect 43250 2970 43340 2990
rect 43250 2930 43270 2970
rect 43320 2930 43340 2970
rect 43250 2920 43340 2930
rect 43250 2890 43300 2920
rect 25790 1820 27370 1840
rect 32190 2850 43300 2890
rect 32190 2800 32230 2850
rect 37050 2800 37090 2850
rect 43450 2800 43490 3050
rect 43660 2970 43750 2990
rect 43660 2930 43680 2970
rect 43730 2930 43750 2970
rect 43660 2920 43750 2930
rect 43690 2890 43750 2920
rect 67680 2890 67720 4880
rect 67770 4800 67860 4820
rect 67770 4760 67790 4800
rect 67840 4790 67860 4800
rect 67840 4760 67890 4790
rect 67770 4750 67890 4760
rect 43690 2850 67720 2890
rect 51390 2800 51430 2850
rect 56250 2800 56290 2850
rect 32190 2780 33770 2800
rect 3270 1680 3310 1820
rect 8970 1680 9010 1820
rect 13490 1690 13580 1710
rect 13490 1680 13510 1690
rect 3270 1650 13510 1680
rect 13560 1650 13580 1690
rect 3270 1640 13580 1650
rect 13490 1560 13580 1580
rect 13490 1550 13510 1560
rect -6400 1520 13510 1550
rect 13560 1520 13580 1560
rect -6400 1510 13580 1520
rect 12920 1440 13010 1460
rect 12920 1430 12940 1440
rect 11330 1400 12940 1430
rect 12990 1430 13010 1440
rect 13490 1440 13580 1460
rect 13490 1430 13510 1440
rect 12990 1400 13510 1430
rect 13560 1400 13580 1440
rect 11330 1390 13580 1400
rect 0 1330 90 1350
rect 0 1290 20 1330
rect 70 1320 90 1330
rect 4860 1330 4950 1350
rect 4860 1320 4880 1330
rect 70 1290 4880 1320
rect 4930 1320 4950 1330
rect 8060 1330 8150 1350
rect 8060 1320 8080 1330
rect 4930 1290 8080 1320
rect 8130 1320 8150 1330
rect 11180 1330 11270 1350
rect 11180 1320 11200 1330
rect 8130 1290 11200 1320
rect 11250 1290 11270 1330
rect 0 1280 11270 1290
rect 9670 1190 9710 1280
rect 11330 1190 11370 1390
rect 11480 1330 11570 1350
rect 11480 1290 11500 1330
rect 11550 1320 11570 1330
rect 13680 1320 13720 1820
rect 13860 1690 13950 1710
rect 13860 1650 13880 1690
rect 13930 1680 13950 1690
rect 18310 1680 18350 1820
rect 24010 1680 24050 1820
rect 13930 1650 24050 1680
rect 13860 1640 24050 1650
rect 32190 1640 32210 2780
rect 33750 1640 33770 2780
rect 13860 1560 13950 1580
rect 13860 1520 13880 1560
rect 13930 1550 13950 1560
rect 18100 1560 18190 1580
rect 18100 1550 18120 1560
rect 13930 1520 18120 1550
rect 18170 1520 18190 1560
rect 13860 1510 18190 1520
rect 13860 1440 13950 1460
rect 13860 1400 13880 1440
rect 13930 1430 13950 1440
rect 18310 1430 18350 1640
rect 32190 1620 33770 1640
rect 35390 2780 36970 2800
rect 35390 1640 35410 2780
rect 36950 1640 36970 2780
rect 35390 1620 36970 1640
rect 37050 2780 38630 2800
rect 37050 1640 37070 2780
rect 38610 1640 38630 2780
rect 37050 1620 38630 1640
rect 40250 2780 41830 2800
rect 40250 1640 40270 2780
rect 41810 1640 41830 2780
rect 40250 1620 41830 1640
rect 43450 2780 45030 2800
rect 43450 1640 43470 2780
rect 45010 1640 45030 2780
rect 43450 1620 45030 1640
rect 46650 2780 48230 2800
rect 46650 1640 46670 2780
rect 48210 1640 48230 2780
rect 46650 1620 48230 1640
rect 49850 2780 51430 2800
rect 49850 1640 49870 2780
rect 51410 1640 51430 2780
rect 49850 1620 51430 1640
rect 51510 2780 53090 2800
rect 51510 1640 51530 2780
rect 53070 1640 53090 2780
rect 51510 1620 53090 1640
rect 54710 2780 56290 2800
rect 54710 1640 54730 2780
rect 56270 1640 56290 2780
rect 54710 1620 56290 1640
rect 57910 2780 61090 2800
rect 57910 1640 57930 2780
rect 59470 1640 59530 2780
rect 61070 1640 61090 2780
rect 57910 1620 61090 1640
rect 57910 1580 57950 1620
rect 18430 1560 18520 1580
rect 18430 1520 18450 1560
rect 18500 1550 18520 1560
rect 33780 1570 33870 1580
rect 33780 1550 33800 1570
rect 18500 1530 33800 1550
rect 33850 1550 33870 1570
rect 38640 1570 38730 1580
rect 38640 1550 38660 1570
rect 33850 1530 38660 1550
rect 38710 1550 38730 1570
rect 41840 1570 41930 1580
rect 41840 1550 41860 1570
rect 38710 1530 41860 1550
rect 41910 1550 41930 1570
rect 46550 1570 46640 1580
rect 46550 1550 46570 1570
rect 41910 1530 46570 1550
rect 46620 1550 46640 1570
rect 49750 1570 49840 1580
rect 49750 1550 49770 1570
rect 46620 1530 49770 1550
rect 49820 1550 49840 1570
rect 54610 1570 54700 1580
rect 54610 1550 54630 1570
rect 49820 1530 54630 1550
rect 54680 1530 54700 1570
rect 18500 1520 54700 1530
rect 18430 1510 54700 1520
rect 57760 1570 57950 1580
rect 57760 1530 57780 1570
rect 57830 1540 57950 1570
rect 57830 1530 57850 1540
rect 57760 1510 57850 1530
rect 20980 1440 21070 1460
rect 20980 1430 21000 1440
rect 13930 1400 21000 1430
rect 21050 1430 21070 1440
rect 38490 1440 38580 1460
rect 38490 1430 38510 1440
rect 21050 1400 38510 1430
rect 38560 1430 38580 1440
rect 46550 1440 46640 1460
rect 46550 1430 46570 1440
rect 38560 1400 46570 1430
rect 46620 1430 46640 1440
rect 46620 1400 67960 1430
rect 13860 1390 67960 1400
rect 16120 1330 16210 1350
rect 16120 1320 16140 1330
rect 11550 1290 16140 1320
rect 16190 1320 16210 1330
rect 19240 1330 19330 1350
rect 19240 1320 19260 1330
rect 16190 1290 19260 1320
rect 19310 1290 19330 1330
rect 11480 1280 19330 1290
rect 17730 1190 17770 1280
rect 19390 1190 19430 1390
rect 19540 1330 19630 1350
rect 19540 1290 19560 1330
rect 19610 1320 19630 1330
rect 24180 1330 24270 1350
rect 24180 1320 24200 1330
rect 19610 1290 24200 1320
rect 24250 1320 24270 1330
rect 27380 1330 27470 1350
rect 27380 1320 27400 1330
rect 24250 1290 27400 1320
rect 27450 1320 27470 1330
rect 32090 1330 32180 1350
rect 32090 1320 32110 1330
rect 27450 1290 32110 1320
rect 32160 1320 32180 1330
rect 35290 1330 35380 1350
rect 35290 1320 35310 1330
rect 32160 1290 35310 1320
rect 35360 1320 35380 1330
rect 39930 1330 40020 1350
rect 39930 1320 39950 1330
rect 35360 1290 39950 1320
rect 40000 1290 40020 1330
rect 19540 1280 40020 1290
rect 25790 1190 25830 1280
rect 33730 1190 33770 1280
rect 40130 1190 40170 1390
rect 40230 1330 40320 1350
rect 40230 1290 40250 1330
rect 40300 1320 40320 1330
rect 43350 1330 43440 1350
rect 43350 1320 43370 1330
rect 40300 1290 43370 1320
rect 43420 1320 43440 1330
rect 47990 1330 48080 1350
rect 47990 1320 48010 1330
rect 43420 1290 48010 1320
rect 48060 1290 48080 1330
rect 40230 1280 48080 1290
rect 41790 1190 41830 1280
rect 48190 1190 48230 1390
rect 48290 1330 48380 1350
rect 48290 1290 48310 1330
rect 48360 1320 48380 1330
rect 51410 1330 51500 1350
rect 51410 1320 51430 1330
rect 48360 1290 51430 1320
rect 51480 1320 51500 1330
rect 54610 1330 54700 1350
rect 54610 1320 54630 1330
rect 51480 1290 54630 1320
rect 54680 1320 54700 1330
rect 59470 1330 59560 1350
rect 59470 1320 59490 1330
rect 54680 1290 59490 1320
rect 59540 1290 59560 1330
rect 48290 1280 59560 1290
rect 49850 1190 49890 1280
rect -6390 1170 -3210 1190
rect -6390 30 -6370 1170
rect -4830 30 -4770 1170
rect -3230 30 -3210 1170
rect -6390 10 -3210 30
rect -1590 1170 -10 1190
rect -1590 30 -1570 1170
rect -30 30 -10 1170
rect -1590 10 -10 30
rect 1610 1170 3190 1190
rect 1610 30 1630 1170
rect 3170 30 3190 1170
rect 1610 10 3190 30
rect 3270 1170 4850 1190
rect 3270 30 3290 1170
rect 4830 30 4850 1170
rect 3270 10 4850 30
rect 6470 1170 8050 1190
rect 6470 30 6490 1170
rect 8030 30 8050 1170
rect 6470 10 8050 30
rect 9670 1170 11250 1190
rect 9670 30 9690 1170
rect 11230 30 11250 1170
rect 9670 10 11250 30
rect 11330 1170 12910 1190
rect 11330 30 11350 1170
rect 12890 30 12910 1170
rect 11330 10 12910 30
rect 14530 1170 16110 1190
rect 14530 30 14550 1170
rect 16090 30 16110 1170
rect 14530 10 16110 30
rect 17730 1170 19310 1190
rect 17730 30 17750 1170
rect 19290 30 19310 1170
rect 17730 10 19310 30
rect 19390 1170 20970 1190
rect 19390 30 19410 1170
rect 20950 30 20970 1170
rect 19390 10 20970 30
rect 22590 1170 24170 1190
rect 22590 30 22610 1170
rect 24150 30 24170 1170
rect 22590 10 24170 30
rect 25790 1170 27370 1190
rect 25790 30 25810 1170
rect 27350 30 27370 1170
rect 25790 10 27370 30
rect 28990 1170 30570 1190
rect 28990 30 29010 1170
rect 30550 30 30570 1170
rect 28990 10 30570 30
rect 32190 1170 33770 1190
rect 32190 30 32210 1170
rect 33750 30 33770 1170
rect 32190 10 33770 30
rect 35390 1170 36970 1190
rect 35390 30 35410 1170
rect 36950 30 36970 1170
rect 35390 10 36970 30
rect 38590 1170 40170 1190
rect 38590 30 38610 1170
rect 40150 30 40170 1170
rect 38590 10 40170 30
rect 40250 1170 41830 1190
rect 40250 30 40270 1170
rect 41810 30 41830 1170
rect 40250 10 41830 30
rect 43450 1170 45030 1190
rect 43450 30 43470 1170
rect 45010 30 45030 1170
rect 43450 10 45030 30
rect 46650 1170 48230 1190
rect 46650 30 46670 1170
rect 48210 30 48230 1170
rect 46650 10 48230 30
rect 48310 1170 49890 1190
rect 48310 30 48330 1170
rect 49870 30 49890 1170
rect 48310 10 49890 30
rect 51510 1170 53090 1190
rect 51510 30 51530 1170
rect 53070 30 53090 1170
rect 51510 10 53090 30
rect 54710 1170 56290 1190
rect 54710 30 54730 1170
rect 56270 30 56290 1170
rect 54710 10 56290 30
rect 56370 1170 57950 1190
rect 56370 30 56390 1170
rect 57930 30 57950 1170
rect 56370 10 57950 30
rect 59570 1170 61150 1190
rect 59570 30 59590 1170
rect 61130 30 61150 1170
rect 59570 10 61150 30
rect 62770 1170 65950 1190
rect 62770 30 62790 1170
rect 64330 30 64390 1170
rect 65930 30 65950 1170
rect 62770 10 65950 30
rect -3250 -30 -3210 10
rect 1610 -30 1650 10
rect 6470 -30 6510 10
rect 14530 -30 14570 10
rect 22590 -30 22630 10
rect 28990 -30 29030 10
rect 36930 -30 36970 10
rect 44990 -30 45030 10
rect 53050 -30 53090 10
rect 57910 -30 57950 10
rect 62770 -30 62810 10
rect -3250 -40 -3110 -30
rect -3250 -70 -3180 -40
rect -3200 -80 -3180 -70
rect -3130 -80 -3110 -40
rect 1610 -70 57950 -30
rect 62670 -40 62810 -30
rect -3200 -100 -3110 -80
rect 62670 -80 62690 -40
rect 62740 -70 62810 -40
rect 62740 -80 62760 -70
rect 62670 -100 62760 -80
<< viali >>
rect -4830 3380 -3290 4520
rect -3230 3380 -1690 4520
rect -30 3380 1510 4520
rect 4830 3380 6370 4520
rect 56270 3380 57810 4520
rect 61130 3380 62670 4520
rect 64330 3380 65870 4520
rect 65930 3380 67470 4520
rect -4830 1840 -3290 2980
rect -3230 1840 -1690 2980
rect -30 1840 1510 2980
rect 4830 1840 6370 2980
rect 9690 1840 11230 2980
rect 16090 1840 17630 2980
rect 20950 1840 22490 2980
rect 25810 1840 27350 2980
rect 35410 1640 36950 2780
rect 40270 1640 41810 2780
rect 46670 1640 48210 2780
rect 51530 1640 53070 2780
rect 57930 1640 59470 2780
rect 59530 1640 61070 2780
rect -6370 30 -4830 1170
rect -4770 30 -3230 1170
rect -1570 30 -30 1170
rect 3290 30 4830 1170
rect 54730 30 56270 1170
rect 59590 30 61130 1170
rect 62790 30 64330 1170
rect 64390 30 65930 1170
<< metal1 >>
rect -4920 4520 67560 4550
rect -4920 3380 -4830 4520
rect -3290 3380 -3230 4520
rect -1690 3380 -30 4520
rect 1510 3380 4830 4520
rect 6370 3380 56270 4520
rect 57810 3380 61130 4520
rect 62670 3380 64330 4520
rect 65870 3380 65930 4520
rect 67470 3380 67560 4520
rect -4920 3350 67560 3380
rect -4920 2980 27450 3350
rect 35190 3280 67560 3350
rect -4920 1840 -4830 2980
rect -3290 1840 -3230 2980
rect -1690 1840 -30 2980
rect 1510 1840 4830 2980
rect 6370 1840 9690 2980
rect 11230 1840 16090 2980
rect 17630 1840 20950 2980
rect 22490 1840 25810 2980
rect 27350 1840 27450 2980
rect -4920 1810 27450 1840
rect 32180 2780 61100 2810
rect 32180 1640 35410 2780
rect 36950 1640 40270 2780
rect 41810 1640 46670 2780
rect 48210 1640 51530 2780
rect 53070 1640 57930 2780
rect 59470 1640 59530 2780
rect 61070 1640 61100 2780
rect 32180 1200 61100 1640
rect -6400 1170 65960 1200
rect -6400 30 -6370 1170
rect -4830 30 -4770 1170
rect -3230 30 -1570 1170
rect -30 30 3290 1170
rect 4830 30 54730 1170
rect 56270 30 59590 1170
rect 61130 30 62790 1170
rect 64330 30 64390 1170
rect 65930 30 65960 1170
rect -6400 0 65960 30
<< labels >>
rlabel locali -6460 3230 -6460 3230 7 Vbp
port 1 w
rlabel locali -6400 1530 -6400 1530 7 Vbn
port 2 w
rlabel locali 67890 4900 67890 4900 3 Vcp
port 3 e
rlabel locali 67960 1410 67960 1410 3 Vcn
port 4 e
rlabel metal1 -6400 1190 -6400 1190 7 VN
port 5 w
rlabel metal1 -4920 1820 -4920 1820 7 VP
port 6 w
<< end >>
