magic
tech sky130A
timestamp 1700326392
<< poly >>
rect 37453 7303 37932 7326
rect 35546 5442 35804 5465
rect 37453 5442 37513 7303
rect 37750 6480 37825 6500
rect 37750 6440 37765 6480
rect 37810 6465 37825 6480
rect 37810 6440 37925 6465
rect 37750 6435 37925 6440
rect 37750 6425 37825 6435
rect 35546 5398 37513 5442
rect 10741 5331 10987 5376
rect 10741 5190 10786 5331
rect 10934 5190 10987 5331
rect 35546 5256 35595 5398
rect 35748 5382 37513 5398
rect 35748 5256 35804 5382
rect 37453 5375 37513 5382
rect 35546 5219 35804 5256
rect 10741 5131 10987 5190
rect 10794 4682 10909 5131
rect 37496 3691 37575 3709
rect 36637 3689 36747 3691
rect 37496 3689 37514 3691
rect 36637 3670 37514 3689
rect 36637 3607 36659 3670
rect 36718 3658 37514 3670
rect 36718 3607 36747 3658
rect 37496 3656 37514 3658
rect 37553 3656 37575 3691
rect 37496 3636 37575 3656
rect 36637 3581 36747 3607
rect 37685 3600 37760 3620
rect 37685 3560 37700 3600
rect 37740 3595 37760 3600
rect 37740 3565 37925 3595
rect 37740 3560 37760 3565
rect 37685 3545 37760 3560
rect -489 3294 -361 3318
rect -489 3212 -465 3294
rect -387 3283 -361 3294
rect -114 3288 7 3312
rect -114 3283 -92 3288
rect -387 3239 -92 3283
rect -387 3212 -361 3239
rect -489 3191 -361 3212
rect -114 3217 -92 3239
rect -13 3217 7 3288
rect -114 3189 7 3217
rect 36822 2892 36934 2915
rect 36822 2824 36843 2892
rect 36905 2880 36934 2892
rect 36905 2849 37920 2880
rect 36905 2824 36934 2849
rect 36822 2803 36934 2824
rect -363 1704 -256 1725
rect -363 1701 -14 1704
rect -363 1643 -337 1701
rect -282 1664 -14 1701
rect -282 1643 -256 1664
rect -363 1613 -256 1643
<< polycont >>
rect 37765 6440 37810 6480
rect 10786 5190 10934 5331
rect 35595 5256 35748 5398
rect 36659 3607 36718 3670
rect 37514 3656 37553 3691
rect 37700 3560 37740 3600
rect -465 3212 -387 3294
rect -92 3217 -13 3288
rect 36843 2824 36905 2892
rect -337 1643 -282 1701
<< locali >>
rect 36965 8670 37410 8690
rect -437 7832 -62 7858
rect -437 3318 -414 7832
rect 37375 7070 37410 8670
rect 37375 7050 37810 7070
rect -338 7005 -89 7006
rect -342 6985 -89 7005
rect -489 3294 -361 3318
rect -489 3212 -465 3294
rect -387 3212 -361 3294
rect -489 3191 -361 3212
rect -342 1725 -316 6985
rect 35546 5398 35804 5465
rect 10741 5331 10987 5376
rect 10741 5190 10786 5331
rect 10934 5190 10987 5331
rect 35546 5256 35595 5398
rect 35748 5395 35804 5398
rect 35546 5253 35597 5256
rect 35750 5253 35804 5395
rect 35546 5219 35804 5253
rect 10741 5131 10987 5190
rect -216 4930 227 4980
rect -363 1701 -256 1725
rect -363 1643 -337 1701
rect -282 1643 -256 1701
rect -363 1613 -256 1643
rect -213 1190 -174 4930
rect 36637 3670 36747 3691
rect 36637 3607 36659 3670
rect 36718 3607 36747 3670
rect 36637 3581 36747 3607
rect -63 3312 -6 3382
rect -114 3288 7 3312
rect -114 3217 -92 3288
rect -13 3217 7 3288
rect -114 3189 7 3217
rect 36651 1358 36684 3581
rect 37030 3580 37065 6945
rect 37770 6500 37810 7050
rect 37750 6480 37825 6500
rect 37750 6440 37765 6480
rect 37810 6440 37825 6480
rect 37750 6425 37825 6440
rect 37557 3709 38008 3748
rect 37496 3691 38008 3709
rect 37496 3656 37514 3691
rect 37553 3685 38008 3691
rect 37553 3656 37575 3685
rect 37496 3636 37575 3656
rect 37685 3600 37760 3620
rect 37685 3580 37700 3600
rect 37030 3560 37700 3580
rect 37740 3560 37760 3600
rect 37030 3550 37760 3560
rect 37685 3545 37760 3550
rect 36822 2892 36934 2915
rect 36822 2824 36843 2892
rect 36905 2824 36934 2892
rect 36822 2803 36934 2824
rect 36831 1423 36869 2803
rect 58618 1423 58639 1427
rect 36831 1398 58639 1423
rect 58543 1358 58566 1359
rect 36651 1329 58566 1358
rect -213 1167 -35 1190
rect 58543 495 58566 1329
rect 58453 476 58566 495
rect 58543 475 58566 476
rect 58618 458 58639 1398
rect 58500 437 58640 458
rect 7020 40 7040 360
rect 7875 40 7895 375
rect 7020 20 7315 40
rect 7450 20 7895 40
rect 14245 40 14265 385
rect 15105 40 15125 360
rect 21475 40 21495 365
rect 22335 40 22355 360
rect 14245 20 14560 40
rect 14695 20 15130 40
rect 21475 20 21855 40
rect 21915 20 22355 40
rect 28705 40 28725 380
rect 29565 40 29585 365
rect 28705 20 29045 40
rect 29180 20 29585 40
rect 35935 40 35955 370
rect 36795 40 36815 365
rect 35935 20 36315 40
rect 36410 20 36815 40
rect 43165 40 43185 360
rect 44025 40 44045 365
rect 43165 20 43575 40
rect 43680 20 44045 40
rect 50395 40 50415 360
rect 51255 40 51275 360
rect 50395 20 50770 40
rect 50905 20 51275 40
<< viali >>
rect 10786 5190 10934 5331
rect 35597 5256 35748 5395
rect 35748 5256 35750 5395
rect 35597 5253 35750 5256
<< metal1 >>
rect -335 8715 -255 8730
rect -335 7115 865 8715
rect -335 4960 -255 7115
rect 35546 5395 35804 5465
rect 10738 5369 10981 5380
rect 35546 5369 35597 5395
rect 10734 5331 35597 5369
rect 10734 5294 10786 5331
rect 10738 5190 10786 5294
rect 10934 5294 35597 5331
rect 10934 5190 10981 5294
rect 35546 5253 35597 5294
rect 35750 5253 35804 5395
rect 35546 5219 35804 5253
rect 10738 5126 10981 5190
rect -335 3480 250 4960
rect -320 1125 -215 3480
rect -65 1290 100 1830
rect -320 1050 105 1125
rect 58480 305 58700 310
rect 7230 220 58700 305
rect 7230 215 58360 220
rect 7020 60 58525 145
rect 7020 55 8565 60
use cascode_voltage_gen  cascode_voltage_gen_0
timestamp 1700317815
transform 1 0 3065 0 1 6230
box -3230 -195 33980 2525
use curgen_1  curgen_1_0
timestamp 1700276151
transform 1 0 3462 0 1 3489
box -3520 -1825 31825 1530
use fvf  fvf_0
timestamp 1700318556
transform 1 0 39675 0 1 430
box -1790 1030 18445 8265
use inverter  inverter_0
timestamp 1700276902
transform 1 0 50980 0 1 145
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1700276902
transform 1 0 7480 0 1 145
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1700276902
transform 1 0 14730 0 1 145
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1700276902
transform 1 0 21980 0 1 145
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1700276902
transform 1 0 29230 0 1 145
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1700276902
transform 1 0 36480 0 1 145
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1700276902
transform 1 0 43730 0 1 145
box -240 -145 -30 185
use ladder  ladder_0
timestamp 1700322215
transform 1 0 10310 0 1 985
box -10460 -640 48280 315
<< end >>
