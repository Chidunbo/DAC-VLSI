magic
tech sky130A
timestamp 1700364827
<< poly >>
rect 36860 7300 38075 7325
rect -695 7085 -625 7100
rect -695 7050 -680 7085
rect -640 7080 -625 7085
rect -140 7090 -70 7105
rect -140 7080 -125 7090
rect -640 7055 -125 7080
rect -85 7055 -70 7090
rect -640 7050 -625 7055
rect -695 7035 -625 7050
rect -140 7040 -70 7055
rect 36690 6520 36750 6525
rect 36860 6520 36910 7300
rect 36690 6465 36910 6520
rect 37525 6485 37600 6500
rect 36690 5740 36750 6465
rect 37525 6440 37540 6485
rect 37585 6465 37600 6485
rect 37585 6440 37905 6465
rect 37525 6435 37905 6440
rect 37525 6425 37600 6435
rect 36465 5675 36770 5740
rect 36465 5505 36540 5675
rect 36715 5505 36770 5675
rect 36465 5445 36770 5505
rect 58300 5120 58455 5155
rect 58300 5095 58335 5120
rect 58050 5065 58335 5095
rect 58300 5040 58335 5065
rect 58425 5040 58455 5120
rect 58300 5000 58455 5040
rect 36970 3615 37080 3650
rect 36970 3555 36995 3615
rect 37055 3595 37080 3615
rect 37055 3565 37965 3595
rect 37055 3555 37080 3565
rect 36970 3535 37080 3555
rect -480 3310 -320 3340
rect -480 3215 -445 3310
rect -350 3280 -320 3310
rect -90 3310 65 3335
rect -90 3280 -60 3310
rect -350 3225 -60 3280
rect -350 3215 -320 3225
rect -480 3195 -320 3215
rect -90 3220 -60 3225
rect 30 3220 65 3310
rect -90 3195 65 3220
rect 37615 2905 37730 2935
rect 37615 2845 37640 2905
rect 37705 2880 37730 2905
rect 37705 2850 37960 2880
rect 37705 2845 37730 2850
rect 37615 2820 37730 2845
rect -680 1730 -585 1745
rect -680 1680 -660 1730
rect -605 1705 -585 1730
rect -605 1680 60 1705
rect -680 1665 60 1680
rect -680 1650 -585 1665
<< polycont >>
rect -680 7050 -640 7085
rect -125 7055 -85 7090
rect 37540 6440 37585 6485
rect 36540 5505 36715 5675
rect 58335 5040 58425 5120
rect 36995 3555 37055 3615
rect -445 3215 -350 3310
rect -60 3220 30 3310
rect 37640 2845 37705 2905
rect -660 1680 -605 1730
<< locali >>
rect 36970 8670 37545 8690
rect -465 7855 -430 7860
rect -465 7835 -75 7855
rect -695 7085 -625 7100
rect -695 7050 -680 7085
rect -640 7050 -625 7085
rect -695 7035 -625 7050
rect -680 1745 -660 7035
rect -465 5525 -430 7835
rect -140 7090 -70 7105
rect -140 7055 -125 7090
rect -85 7055 -70 7090
rect -140 7040 -70 7055
rect -135 6985 -105 7040
rect 36475 5675 36775 5740
rect -230 5555 -90 5580
rect -230 5525 -210 5555
rect -465 5470 -210 5525
rect -120 5470 -90 5555
rect -465 3340 -430 5470
rect -230 5440 -90 5470
rect 36475 5505 36540 5675
rect 36715 5505 36775 5675
rect 36475 5450 36775 5505
rect -275 4925 110 4970
rect -480 3310 -320 3340
rect -480 3215 -445 3310
rect -350 3215 -320 3310
rect -480 3195 -320 3215
rect -680 1730 -585 1745
rect -680 1680 -660 1730
rect -605 1680 -585 1730
rect -680 1650 -585 1680
rect -275 1190 -200 4925
rect 36965 3650 37020 6945
rect 37525 6500 37545 8670
rect 37525 6485 37600 6500
rect 37525 6440 37540 6485
rect 37585 6440 37600 6485
rect 37525 6425 37600 6440
rect 37525 6420 37545 6425
rect 58300 5120 58455 5155
rect 58300 5040 58335 5120
rect 58425 5040 58455 5120
rect 58300 5000 58455 5040
rect 37240 3690 37990 3750
rect 36965 3615 37080 3650
rect 36965 3585 36995 3615
rect 36970 3555 36995 3585
rect 37055 3555 37080 3615
rect 36970 3535 37080 3555
rect -60 3335 15 3395
rect -90 3310 65 3335
rect -90 3220 -60 3310
rect 30 3220 65 3310
rect -90 3195 65 3220
rect 37240 1865 37305 3690
rect 37615 2905 37730 2935
rect 37615 2845 37640 2905
rect 37705 2845 37730 2905
rect 37615 2820 37730 2845
rect 37245 1340 37305 1865
rect 37680 1430 37715 2820
rect 37680 1395 58745 1430
rect 37685 1385 58745 1395
rect 58635 1380 58745 1385
rect 37245 1300 58640 1340
rect -275 1170 -70 1190
rect 58615 495 58640 1300
rect 58510 475 58640 495
rect 58710 455 58745 1380
rect 58495 435 58745 455
rect 7014 40 7035 382
rect 7876 40 7897 356
rect 14245 40 14266 352
rect 7013 19 7286 40
rect 7434 19 7898 40
rect 14245 17 14525 40
rect 15106 39 15127 370
rect 21475 41 21495 366
rect 22335 41 22357 362
rect 14659 18 15147 39
rect 21475 18 21774 41
rect 22220 40 22357 41
rect 21935 20 22357 40
rect 28705 39 28727 381
rect 29564 43 29586 354
rect 29483 41 29601 43
rect 22220 19 22353 20
rect 28702 18 29025 39
rect 29190 20 29601 41
rect 35935 40 35955 360
rect 36795 40 36815 360
rect 35935 20 36315 40
rect 36435 20 36815 40
rect 43165 40 43185 360
rect 44025 40 44045 360
rect 50395 40 50415 355
rect 51255 40 51275 360
rect 43165 20 43545 40
rect 43685 20 44065 40
rect 50395 20 50800 40
rect 50395 15 50415 20
rect 50930 20 51290 40
<< viali >>
rect -210 5470 -120 5555
rect 36540 5510 36715 5675
rect 58335 5040 58425 5120
rect 7345 10 7365 30
rect 14595 10 14615 30
rect 21845 10 21865 30
rect 29095 10 29115 30
rect 36345 10 36365 30
rect 43595 10 43615 30
rect 50845 10 50865 30
<< metal1 >>
rect -415 8670 1280 8685
rect -440 7135 1280 8670
rect 36655 7860 38410 8700
rect -440 4950 -310 7135
rect 37175 6395 37330 6410
rect 35980 6255 37330 6395
rect 36475 5675 36775 5740
rect -240 5555 -40 5610
rect -240 5470 -210 5555
rect -120 5550 -40 5555
rect 36475 5550 36540 5675
rect -120 5510 36540 5550
rect 36715 5510 36775 5675
rect -120 5470 36775 5510
rect -240 5405 -40 5470
rect 36475 5450 36775 5470
rect -440 4640 105 4950
rect -425 3475 105 4640
rect 37175 4125 37330 6255
rect 58295 5120 58460 5160
rect 58295 5040 58335 5120
rect 58425 5080 58460 5120
rect 58425 5040 58820 5080
rect 58295 5015 58820 5040
rect 58295 5005 58460 5015
rect 37175 3950 37945 4125
rect -425 1125 -325 3475
rect 28685 1275 29205 1805
rect 35245 1745 38215 3115
rect 58505 1175 58825 1310
rect -425 1045 235 1125
rect -425 330 -325 1045
rect -425 325 105 330
rect -425 210 58615 325
rect -425 205 105 210
rect 58725 155 58820 1175
rect 58570 150 58820 155
rect -130 75 58820 150
rect 7335 30 7375 40
rect 7335 10 7345 30
rect 7365 10 7375 30
rect 7335 -65 7375 10
rect 14585 30 14625 40
rect 14585 10 14595 30
rect 14615 10 14625 30
rect 14585 -65 14625 10
rect 21835 30 21875 40
rect 21835 10 21845 30
rect 21865 10 21875 30
rect 21835 -65 21875 10
rect 29085 30 29125 40
rect 29085 10 29095 30
rect 29115 10 29125 30
rect 29085 -65 29125 10
rect 36335 30 36375 40
rect 36335 10 36345 30
rect 36365 10 36375 30
rect 36335 -65 36375 10
rect 43585 30 43625 40
rect 43585 10 43595 30
rect 43615 10 43625 30
rect 43585 -65 43625 10
rect 50835 30 50875 40
rect 50835 10 50845 30
rect 50865 10 50875 30
rect 50835 -65 50875 10
use FVF_lds  FVF_lds_0
timestamp 1700362378
transform 1 0 39675 0 1 430
box -1790 1030 18445 8265
use inverter  inverter_0
timestamp 1700276902
transform 1 0 50980 0 1 145
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1700276902
transform 1 0 7480 0 1 145
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1700276902
transform 1 0 14730 0 1 145
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1700276902
transform 1 0 21980 0 1 145
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1700276902
transform 1 0 29230 0 1 145
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1700276902
transform 1 0 36480 0 1 145
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1700276902
transform 1 0 43730 0 1 145
box -240 -145 -30 185
use lds-curgen-j1  lds-curgen-j1_0
timestamp 1700276151
transform 1 0 3462 0 1 3489
box -3520 -1825 31825 1530
use lds-ladder  lds-ladder_0
timestamp 1700322215
transform 1 0 10310 0 1 985
box -10460 -640 48280 315
use VGen  VGen_0
timestamp 1700345324
transform 1 0 3065 0 1 6230
box -3230 -105 33980 2525
<< labels >>
rlabel metal1 58820 5050 58820 5050 3 Ifout
rlabel metal1 -130 90 -130 90 7 VN
rlabel metal1 -425 265 -425 265 7 VP
rlabel metal1 7354 -65 7354 -65 5 Vin6
rlabel metal1 14605 -65 14605 -65 5 Vin5
rlabel metal1 21853 -65 21853 -65 5 Vin4
rlabel metal1 29105 -65 29105 -65 5 Vin3
rlabel metal1 36352 -65 36352 -65 5 Vin2
rlabel metal1 43606 -65 43606 -65 5 Vin1
rlabel metal1 50855 -65 50855 -65 5 Vin0
<< end >>
