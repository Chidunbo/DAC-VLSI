magic
tech sky130A
timestamp 1700276902
<< nwell >>
rect 2385 8585 2540 8640
rect 4885 8585 5040 8640
rect 7385 8585 7540 8640
rect 9885 8585 10040 8640
rect 11735 8585 11890 8640
rect 13885 8585 14040 8640
rect 15785 8585 15940 8640
rect 17885 8585 18040 8640
rect 19935 8585 20090 8640
rect 21885 8585 22040 8640
rect 23885 8585 24040 8640
rect 25885 8585 26040 8640
rect 27885 8585 28040 8640
rect 29885 8585 30040 8640
rect 31885 8585 32040 8640
rect 33915 8555 34010 8575
<< psubdiff >>
rect 17720 7725 17875 7740
rect 17720 7705 17745 7725
rect 17850 7705 17875 7725
rect 17720 7685 17875 7705
rect 20720 7725 20875 7740
rect 20720 7705 20745 7725
rect 20850 7705 20875 7725
rect 20720 7685 20875 7705
rect 23720 7725 23875 7740
rect 23720 7705 23745 7725
rect 23850 7705 23875 7725
rect 23720 7685 23875 7705
rect 26720 7725 26875 7740
rect 26720 7705 26745 7725
rect 26850 7705 26875 7725
rect 26720 7685 26875 7705
rect 28720 7725 28875 7740
rect 28720 7705 28745 7725
rect 28850 7705 28875 7725
rect 28720 7685 28875 7705
rect 30720 7725 30875 7740
rect 30720 7705 30745 7725
rect 30850 7705 30875 7725
rect 30720 7685 30875 7705
rect 3335 6105 3490 6120
rect 3335 6085 3365 6105
rect 3460 6085 3490 6105
rect 3335 6065 3490 6085
rect 5335 6105 5490 6120
rect 5335 6085 5365 6105
rect 5460 6085 5490 6105
rect 5335 6065 5490 6085
rect 7335 6105 7490 6120
rect 7335 6085 7365 6105
rect 7460 6085 7490 6105
rect 7335 6065 7490 6085
rect 9335 6105 9490 6120
rect 9335 6085 9365 6105
rect 9460 6085 9490 6105
rect 9335 6065 9490 6085
rect 11335 6105 11490 6120
rect 11335 6085 11365 6105
rect 11460 6085 11490 6105
rect 11335 6065 11490 6085
rect 13335 6105 13490 6120
rect 13335 6085 13365 6105
rect 13460 6085 13490 6105
rect 13335 6065 13490 6085
rect 15335 6105 15490 6120
rect 15335 6085 15365 6105
rect 15460 6085 15490 6105
rect 15335 6065 15490 6085
rect 17335 6105 17490 6120
rect 17335 6085 17365 6105
rect 17460 6085 17490 6105
rect 17335 6065 17490 6085
rect 19335 6105 19490 6120
rect 19335 6085 19365 6105
rect 19460 6085 19490 6105
rect 19335 6065 19490 6085
rect 3200 1285 3300 1300
rect 3200 1265 3215 1285
rect 3285 1265 3300 1285
rect 3200 1250 3300 1265
rect 5200 1285 5300 1300
rect 5200 1265 5215 1285
rect 5285 1265 5300 1285
rect 5200 1250 5300 1265
rect 7200 1285 7300 1300
rect 7200 1265 7215 1285
rect 7285 1265 7300 1285
rect 7200 1250 7300 1265
rect 9200 1285 9300 1300
rect 9200 1265 9215 1285
rect 9285 1265 9300 1285
rect 9200 1250 9300 1265
rect 11200 1285 11300 1300
rect 11200 1265 11215 1285
rect 11285 1265 11300 1285
rect 11200 1250 11300 1265
rect 13200 1285 13300 1300
rect 13200 1265 13215 1285
rect 13285 1265 13300 1285
rect 13200 1250 13300 1265
rect 15200 1285 15300 1300
rect 15200 1265 15215 1285
rect 15285 1265 15300 1285
rect 15200 1250 15300 1265
rect 17200 1285 17300 1300
rect 17200 1265 17215 1285
rect 17285 1265 17300 1285
rect 17200 1250 17300 1265
rect 19200 1285 19300 1300
rect 19200 1265 19215 1285
rect 19285 1265 19300 1285
rect 19200 1250 19300 1265
rect 21200 1285 21300 1300
rect 21200 1265 21215 1285
rect 21285 1265 21300 1285
rect 21200 1250 21300 1265
rect 23200 1285 23300 1300
rect 23200 1265 23215 1285
rect 23285 1265 23300 1285
rect 23200 1250 23300 1265
rect 25200 1285 25300 1300
rect 25200 1265 25215 1285
rect 25285 1265 25300 1285
rect 25200 1250 25300 1265
rect 27200 1285 27300 1300
rect 27200 1265 27215 1285
rect 27285 1265 27300 1285
rect 27200 1250 27300 1265
rect 29200 1285 29300 1300
rect 29200 1265 29215 1285
rect 29285 1265 29300 1285
rect 29200 1250 29300 1265
rect 31200 1285 31300 1300
rect 31200 1265 31215 1285
rect 31285 1265 31300 1285
rect 31200 1250 31300 1265
rect 33200 1285 33300 1300
rect 33200 1265 33215 1285
rect 33285 1265 33300 1285
rect 33200 1250 33300 1265
rect 35200 1285 35300 1300
rect 35200 1265 35215 1285
rect 35285 1265 35300 1285
rect 35200 1250 35300 1265
rect 37200 1285 37300 1300
rect 37200 1265 37215 1285
rect 37285 1265 37300 1285
rect 37200 1250 37300 1265
rect 39200 1285 39300 1300
rect 39200 1265 39215 1285
rect 39285 1265 39300 1285
rect 39200 1250 39300 1265
rect 41200 1285 41300 1300
rect 41200 1265 41215 1285
rect 41285 1265 41300 1285
rect 41200 1250 41300 1265
rect 43200 1285 43300 1300
rect 43200 1265 43215 1285
rect 43285 1265 43300 1285
rect 43200 1250 43300 1265
rect 45200 1285 45300 1300
rect 45200 1265 45215 1285
rect 45285 1265 45300 1285
rect 45200 1250 45300 1265
rect 47200 1285 47300 1300
rect 47200 1265 47215 1285
rect 47285 1265 47300 1285
rect 47200 1250 47300 1265
rect 49200 1285 49300 1300
rect 49200 1265 49215 1285
rect 49285 1265 49300 1285
rect 49200 1250 49300 1265
rect 53550 1285 53650 1300
rect 53550 1265 53565 1285
rect 53635 1265 53650 1285
rect 53550 1250 53650 1265
rect 57550 1285 57650 1300
rect 57550 1265 57565 1285
rect 57635 1265 57650 1285
rect 57550 1250 57650 1265
<< nsubdiff >>
rect 2385 8625 2540 8640
rect 2385 8605 2415 8625
rect 2510 8605 2540 8625
rect 2385 8585 2540 8605
rect 4885 8625 5040 8640
rect 4885 8605 4915 8625
rect 5010 8605 5040 8625
rect 4885 8585 5040 8605
rect 7385 8625 7540 8640
rect 7385 8605 7415 8625
rect 7510 8605 7540 8625
rect 7385 8585 7540 8605
rect 9885 8625 10040 8640
rect 9885 8605 9915 8625
rect 10010 8605 10040 8625
rect 9885 8585 10040 8605
rect 11735 8625 11890 8640
rect 11735 8605 11765 8625
rect 11860 8605 11890 8625
rect 11735 8585 11890 8605
rect 13885 8625 14040 8640
rect 13885 8605 13915 8625
rect 14010 8605 14040 8625
rect 13885 8585 14040 8605
rect 15785 8625 15940 8640
rect 15785 8605 15815 8625
rect 15910 8605 15940 8625
rect 15785 8585 15940 8605
rect 17885 8625 18040 8640
rect 17885 8605 17915 8625
rect 18010 8605 18040 8625
rect 17885 8585 18040 8605
rect 19935 8625 20090 8640
rect 19935 8605 19965 8625
rect 20060 8605 20090 8625
rect 19935 8585 20090 8605
rect 21885 8625 22040 8640
rect 21885 8605 21915 8625
rect 22010 8605 22040 8625
rect 21885 8585 22040 8605
rect 23885 8625 24040 8640
rect 23885 8605 23915 8625
rect 24010 8605 24040 8625
rect 23885 8585 24040 8605
rect 25885 8625 26040 8640
rect 25885 8605 25915 8625
rect 26010 8605 26040 8625
rect 25885 8585 26040 8605
rect 27885 8625 28040 8640
rect 27885 8605 27915 8625
rect 28010 8605 28040 8625
rect 27885 8585 28040 8605
rect 29885 8625 30040 8640
rect 29885 8605 29915 8625
rect 30010 8605 30040 8625
rect 29885 8585 30040 8605
rect 31885 8625 32040 8640
rect 31885 8605 31915 8625
rect 32010 8605 32040 8625
rect 31885 8585 32040 8605
rect 33885 8575 34040 8590
rect 33885 8555 33915 8575
rect 34010 8555 34040 8575
rect 33885 8535 34040 8555
<< psubdiffcont >>
rect 17745 7705 17850 7725
rect 20745 7705 20850 7725
rect 23745 7705 23850 7725
rect 26745 7705 26850 7725
rect 28745 7705 28850 7725
rect 30745 7705 30850 7725
rect 3365 6085 3460 6105
rect 5365 6085 5460 6105
rect 7365 6085 7460 6105
rect 9365 6085 9460 6105
rect 11365 6085 11460 6105
rect 13365 6085 13460 6105
rect 15365 6085 15460 6105
rect 17365 6085 17460 6105
rect 19365 6085 19460 6105
rect 3215 1265 3285 1285
rect 5215 1265 5285 1285
rect 7215 1265 7285 1285
rect 9215 1265 9285 1285
rect 11215 1265 11285 1285
rect 13215 1265 13285 1285
rect 15215 1265 15285 1285
rect 17215 1265 17285 1285
rect 19215 1265 19285 1285
rect 21215 1265 21285 1285
rect 23215 1265 23285 1285
rect 25215 1265 25285 1285
rect 27215 1265 27285 1285
rect 29215 1265 29285 1285
rect 31215 1265 31285 1285
rect 33215 1265 33285 1285
rect 35215 1265 35285 1285
rect 37215 1265 37285 1285
rect 39215 1265 39285 1285
rect 41215 1265 41285 1285
rect 43215 1265 43285 1285
rect 45215 1265 45285 1285
rect 47215 1265 47285 1285
rect 49215 1265 49285 1285
rect 53565 1265 53635 1285
rect 57565 1265 57635 1285
<< nsubdiffcont >>
rect 2415 8605 2510 8625
rect 4915 8605 5010 8625
rect 7415 8605 7510 8625
rect 9915 8605 10010 8625
rect 11765 8605 11860 8625
rect 13915 8605 14010 8625
rect 15815 8605 15910 8625
rect 17915 8605 18010 8625
rect 19965 8605 20060 8625
rect 21915 8605 22010 8625
rect 23915 8605 24010 8625
rect 25915 8605 26010 8625
rect 27915 8605 28010 8625
rect 29915 8605 30010 8625
rect 31915 8605 32010 8625
rect 33915 8555 34010 8575
<< poly >>
rect 37750 6480 37825 6500
rect 37750 6440 37765 6480
rect 37810 6465 37825 6480
rect 37810 6440 37925 6465
rect 37750 6435 37925 6440
rect 37750 6425 37825 6435
rect 37685 3600 37760 3620
rect 37685 3560 37700 3600
rect 37740 3595 37760 3600
rect 37740 3565 37925 3595
rect 37740 3560 37760 3565
rect 37685 3545 37760 3560
<< polycont >>
rect 37765 6440 37810 6480
rect 37700 3560 37740 3600
<< locali >>
rect 2400 8625 2525 8630
rect 2400 8605 2415 8625
rect 2510 8605 2525 8625
rect 2400 8595 2525 8605
rect 4900 8625 5025 8630
rect 4900 8605 4915 8625
rect 5010 8605 5025 8625
rect 4900 8595 5025 8605
rect 7400 8625 7525 8630
rect 7400 8605 7415 8625
rect 7510 8605 7525 8625
rect 7400 8595 7525 8605
rect 9900 8625 10025 8630
rect 9900 8605 9915 8625
rect 10010 8605 10025 8625
rect 9900 8595 10025 8605
rect 11750 8625 11875 8630
rect 11750 8605 11765 8625
rect 11860 8605 11875 8625
rect 11750 8595 11875 8605
rect 13900 8625 14025 8630
rect 13900 8605 13915 8625
rect 14010 8605 14025 8625
rect 13900 8595 14025 8605
rect 15800 8625 15925 8630
rect 15800 8605 15815 8625
rect 15910 8605 15925 8625
rect 15800 8595 15925 8605
rect 17900 8625 18025 8630
rect 17900 8605 17915 8625
rect 18010 8605 18025 8625
rect 17900 8595 18025 8605
rect 19950 8625 20075 8630
rect 19950 8605 19965 8625
rect 20060 8605 20075 8625
rect 19950 8595 20075 8605
rect 21900 8625 22025 8630
rect 21900 8605 21915 8625
rect 22010 8605 22025 8625
rect 21900 8595 22025 8605
rect 23900 8625 24025 8630
rect 23900 8605 23915 8625
rect 24010 8605 24025 8625
rect 23900 8595 24025 8605
rect 25900 8625 26025 8630
rect 25900 8605 25915 8625
rect 26010 8605 26025 8625
rect 25900 8595 26025 8605
rect 27900 8625 28025 8630
rect 27900 8605 27915 8625
rect 28010 8605 28025 8625
rect 27900 8595 28025 8605
rect 29900 8625 30025 8630
rect 29900 8605 29915 8625
rect 30010 8605 30025 8625
rect 29900 8595 30025 8605
rect 31900 8625 32025 8630
rect 31900 8605 31915 8625
rect 32010 8605 32025 8625
rect 31900 8595 32025 8605
rect 33900 8575 34025 8580
rect 33900 8555 33915 8575
rect 34010 8555 34025 8575
rect 33900 8545 34025 8555
rect 17730 7725 17865 7730
rect 17730 7705 17745 7725
rect 17850 7705 17865 7725
rect 17730 7695 17865 7705
rect 20730 7725 20865 7730
rect 20730 7705 20745 7725
rect 20850 7705 20865 7725
rect 20730 7695 20865 7705
rect 23730 7725 23865 7730
rect 23730 7705 23745 7725
rect 23850 7705 23865 7725
rect 23730 7695 23865 7705
rect 26730 7725 26865 7730
rect 26730 7705 26745 7725
rect 26850 7705 26865 7725
rect 26730 7695 26865 7705
rect 28730 7725 28865 7730
rect 28730 7705 28745 7725
rect 28850 7705 28865 7725
rect 28730 7695 28865 7705
rect 30730 7725 30865 7730
rect 30730 7705 30745 7725
rect 30850 7705 30865 7725
rect 30730 7695 30865 7705
rect 36905 7070 36925 7685
rect 36905 7050 37810 7070
rect 3350 6105 3475 6110
rect 3350 6085 3365 6105
rect 3460 6085 3475 6105
rect 3350 6075 3475 6085
rect 5350 6105 5475 6110
rect 5350 6085 5365 6105
rect 5460 6085 5475 6105
rect 5350 6075 5475 6085
rect 7350 6105 7475 6110
rect 7350 6085 7365 6105
rect 7460 6085 7475 6105
rect 7350 6075 7475 6085
rect 9350 6105 9475 6110
rect 9350 6085 9365 6105
rect 9460 6085 9475 6105
rect 9350 6075 9475 6085
rect 11350 6105 11475 6110
rect 11350 6085 11365 6105
rect 11460 6085 11475 6105
rect 11350 6075 11475 6085
rect 13350 6105 13475 6110
rect 13350 6085 13365 6105
rect 13460 6085 13475 6105
rect 13350 6075 13475 6085
rect 15350 6105 15475 6110
rect 15350 6085 15365 6105
rect 15460 6085 15475 6105
rect 15350 6075 15475 6085
rect 17350 6105 17475 6110
rect 17350 6085 17365 6105
rect 17460 6085 17475 6105
rect 17350 6075 17475 6085
rect 19350 6105 19475 6110
rect 19350 6085 19365 6105
rect 19460 6085 19475 6105
rect 19350 6075 19475 6085
rect 37030 3580 37065 6945
rect 37770 6500 37810 7050
rect 37750 6480 37825 6500
rect 37750 6440 37765 6480
rect 37810 6440 37825 6480
rect 37750 6425 37825 6440
rect 37685 3600 37760 3620
rect 37685 3580 37700 3600
rect 37030 3560 37700 3580
rect 37740 3560 37760 3600
rect 37030 3550 37760 3560
rect 37685 3545 37760 3550
rect 3205 1285 3295 1295
rect 3205 1265 3215 1285
rect 3285 1265 3295 1285
rect 3205 1255 3295 1265
rect 5205 1285 5295 1295
rect 5205 1265 5215 1285
rect 5285 1265 5295 1285
rect 5205 1255 5295 1265
rect 7205 1285 7295 1295
rect 7205 1265 7215 1285
rect 7285 1265 7295 1285
rect 7205 1255 7295 1265
rect 9205 1285 9295 1295
rect 9205 1265 9215 1285
rect 9285 1265 9295 1285
rect 9205 1255 9295 1265
rect 11205 1285 11295 1295
rect 11205 1265 11215 1285
rect 11285 1265 11295 1285
rect 11205 1255 11295 1265
rect 13205 1285 13295 1295
rect 13205 1265 13215 1285
rect 13285 1265 13295 1285
rect 13205 1255 13295 1265
rect 15205 1285 15295 1295
rect 15205 1265 15215 1285
rect 15285 1265 15295 1285
rect 15205 1255 15295 1265
rect 17205 1285 17295 1295
rect 17205 1265 17215 1285
rect 17285 1265 17295 1285
rect 17205 1255 17295 1265
rect 19205 1285 19295 1295
rect 19205 1265 19215 1285
rect 19285 1265 19295 1285
rect 19205 1255 19295 1265
rect 21205 1285 21295 1295
rect 21205 1265 21215 1285
rect 21285 1265 21295 1285
rect 21205 1255 21295 1265
rect 23205 1285 23295 1295
rect 23205 1265 23215 1285
rect 23285 1265 23295 1285
rect 23205 1255 23295 1265
rect 25205 1285 25295 1295
rect 25205 1265 25215 1285
rect 25285 1265 25295 1285
rect 25205 1255 25295 1265
rect 27205 1285 27295 1295
rect 27205 1265 27215 1285
rect 27285 1265 27295 1285
rect 27205 1255 27295 1265
rect 29205 1285 29295 1295
rect 29205 1265 29215 1285
rect 29285 1265 29295 1285
rect 29205 1255 29295 1265
rect 31205 1285 31295 1295
rect 31205 1265 31215 1285
rect 31285 1265 31295 1285
rect 31205 1255 31295 1265
rect 33205 1285 33295 1295
rect 33205 1265 33215 1285
rect 33285 1265 33295 1285
rect 33205 1255 33295 1265
rect 35205 1285 35295 1295
rect 35205 1265 35215 1285
rect 35285 1265 35295 1285
rect 35205 1255 35295 1265
rect 37205 1285 37295 1295
rect 37205 1265 37215 1285
rect 37285 1265 37295 1285
rect 37205 1255 37295 1265
rect 39205 1285 39295 1295
rect 39205 1265 39215 1285
rect 39285 1265 39295 1285
rect 39205 1255 39295 1265
rect 41205 1285 41295 1295
rect 41205 1265 41215 1285
rect 41285 1265 41295 1285
rect 41205 1255 41295 1265
rect 43205 1285 43295 1295
rect 43205 1265 43215 1285
rect 43285 1265 43295 1285
rect 43205 1255 43295 1265
rect 45205 1285 45295 1295
rect 45205 1265 45215 1285
rect 45285 1265 45295 1285
rect 45205 1255 45295 1265
rect 47205 1285 47295 1295
rect 47205 1265 47215 1285
rect 47285 1265 47295 1285
rect 47205 1255 47295 1265
rect 49205 1285 49295 1295
rect 49205 1265 49215 1285
rect 49285 1265 49295 1285
rect 49205 1255 49295 1265
rect 53555 1285 53645 1295
rect 53555 1265 53565 1285
rect 53635 1265 53645 1285
rect 53555 1255 53645 1265
rect 57555 1285 57645 1295
rect 57555 1265 57565 1285
rect 57635 1265 57645 1285
rect 57555 1255 57645 1265
rect 7015 40 7035 360
rect 7875 40 7895 375
rect 7015 20 7315 40
rect 7450 20 7895 40
rect 14245 40 14265 385
rect 15105 40 15125 360
rect 21475 40 21495 365
rect 22335 40 22355 360
rect 14245 20 14560 40
rect 14695 20 15130 40
rect 21475 20 21855 40
rect 21915 20 22355 40
rect 28705 40 28725 380
rect 29565 40 29585 365
rect 28705 20 29045 40
rect 29180 20 29585 40
rect 35935 40 35955 370
rect 36795 40 36815 365
rect 35935 20 36315 40
rect 36410 20 36815 40
rect 43165 40 43185 360
rect 44025 40 44045 365
rect 43165 20 43575 40
rect 43680 20 44045 40
rect 50395 40 50415 360
rect 51255 40 51275 360
rect 50395 20 50770 40
rect 50905 20 51275 40
<< viali >>
rect 2415 8605 2510 8625
rect 4915 8605 5010 8625
rect 7415 8605 7510 8625
rect 9915 8605 10010 8625
rect 11765 8605 11860 8625
rect 13915 8605 14010 8625
rect 15815 8605 15910 8625
rect 17915 8605 18010 8625
rect 19965 8605 20060 8625
rect 21915 8605 22010 8625
rect 23915 8605 24010 8625
rect 25915 8605 26010 8625
rect 27915 8605 28010 8625
rect 29915 8605 30010 8625
rect 31915 8605 32010 8625
rect 33915 8555 34010 8575
rect 17745 7705 17850 7725
rect 20745 7705 20850 7725
rect 23745 7705 23850 7725
rect 26745 7705 26850 7725
rect 28745 7705 28850 7725
rect 30745 7705 30850 7725
rect 3365 6085 3460 6105
rect 5365 6085 5460 6105
rect 7365 6085 7460 6105
rect 9365 6085 9460 6105
rect 11365 6085 11460 6105
rect 13365 6085 13460 6105
rect 15365 6085 15460 6105
rect 17365 6085 17460 6105
rect 19365 6085 19460 6105
<< metal1 >>
rect 2355 8625 2610 8640
rect 2355 8605 2415 8625
rect 2510 8605 2610 8625
rect 2355 8490 2610 8605
rect 4870 8625 5070 8655
rect 4870 8605 4915 8625
rect 5010 8605 5070 8625
rect 4870 8465 5070 8605
rect 7355 8625 7555 8670
rect 7355 8605 7415 8625
rect 7510 8605 7555 8625
rect 7355 8480 7555 8605
rect 9865 8625 10065 8670
rect 9865 8605 9915 8625
rect 10010 8605 10065 8625
rect 9865 8480 10065 8605
rect 11720 8625 11920 8680
rect 11720 8605 11765 8625
rect 11860 8605 11920 8625
rect 11720 8490 11920 8605
rect 13875 8625 14075 8670
rect 13875 8605 13915 8625
rect 14010 8605 14075 8625
rect 13875 8480 14075 8605
rect 15785 8625 15985 8670
rect 15785 8605 15815 8625
rect 15910 8605 15985 8625
rect 15785 8480 15985 8605
rect 17865 8625 18065 8665
rect 17865 8605 17915 8625
rect 18010 8605 18065 8625
rect 17865 8475 18065 8605
rect 19920 8625 20130 8665
rect 19920 8605 19965 8625
rect 20060 8605 20130 8625
rect 19920 8475 20130 8605
rect 21860 8625 22070 8660
rect 21860 8605 21915 8625
rect 22010 8605 22070 8625
rect 21860 8470 22070 8605
rect 23865 8625 24075 8665
rect 23865 8605 23915 8625
rect 24010 8605 24075 8625
rect 23865 8475 24075 8605
rect 25880 8625 26090 8665
rect 25880 8605 25915 8625
rect 26010 8605 26090 8625
rect 25880 8475 26090 8605
rect 27860 8625 28070 8670
rect 27860 8605 27915 8625
rect 28010 8605 28070 8625
rect 27860 8480 28070 8605
rect 29860 8625 30070 8665
rect 29860 8605 29915 8625
rect 30010 8605 30070 8625
rect 29860 8475 30070 8605
rect 31840 8625 32050 8665
rect 31840 8605 31915 8625
rect 32010 8605 32050 8625
rect 31840 8475 32050 8605
rect 33855 8575 34065 8650
rect 33855 8555 33915 8575
rect 34010 8555 34065 8575
rect 33855 8460 34065 8555
rect 36665 7865 38305 8500
rect 17630 7725 17975 7760
rect 17630 7705 17745 7725
rect 17850 7705 17975 7725
rect 17630 7635 17975 7705
rect 20690 7725 20900 7765
rect 20690 7705 20745 7725
rect 20850 7705 20900 7725
rect 17630 7050 20225 7635
rect 20690 7630 20900 7705
rect 23700 7725 23910 7765
rect 23700 7705 23745 7725
rect 23850 7705 23910 7725
rect 23700 7630 23910 7705
rect 26700 7725 26910 7765
rect 26700 7705 26745 7725
rect 26850 7705 26910 7725
rect 26700 7630 26910 7705
rect 28685 7725 28895 7760
rect 28685 7705 28745 7725
rect 28850 7705 28895 7725
rect 28685 7625 28895 7705
rect 30705 7725 30915 7750
rect 30705 7705 30745 7725
rect 30850 7705 30915 7725
rect 30705 7615 30915 7705
rect 35350 6810 36065 6815
rect 3335 6105 3490 6315
rect 3335 6085 3365 6105
rect 3460 6085 3490 6105
rect 3335 6065 3490 6085
rect 5335 6105 5495 6335
rect 5335 6085 5365 6105
rect 5460 6085 5495 6105
rect 5335 6065 5495 6085
rect 7330 6105 7490 6330
rect 7330 6085 7365 6105
rect 7460 6085 7490 6105
rect 7330 6060 7490 6085
rect 9335 6105 9490 6330
rect 9335 6085 9365 6105
rect 9460 6085 9490 6105
rect 9335 6060 9490 6085
rect 11335 6105 11490 6335
rect 11335 6085 11365 6105
rect 11460 6085 11490 6105
rect 11335 6065 11490 6085
rect 13335 6105 13490 6335
rect 13335 6085 13365 6105
rect 13460 6085 13490 6105
rect 13335 6065 13490 6085
rect 15335 6105 15490 6335
rect 15335 6085 15365 6105
rect 15460 6085 15490 6105
rect 15335 6065 15490 6085
rect 17335 6105 17490 6335
rect 17335 6085 17365 6105
rect 17460 6085 17490 6105
rect 17335 6065 17490 6085
rect 19335 6105 19490 6340
rect 35350 6230 37365 6810
rect 19335 6085 19365 6105
rect 19460 6085 19490 6105
rect 19335 6065 19490 6085
rect 36035 5050 37360 6230
rect 36035 4055 38680 5050
rect 55915 1045 58645 1085
rect -60 145 -5 885
rect 58505 305 58640 1045
rect 7230 215 58640 305
rect 58505 210 58640 215
rect -60 60 58525 145
rect -60 55 8565 60
use cascode_voltage_gen  cascode_voltage_gen_0
timestamp 1700276902
transform 1 0 3065 0 1 6230
box -3230 -50 33980 2525
use fvf  fvf_0
timestamp 1700263747
transform 1 0 39675 0 1 430
box -1790 1030 18445 8265
use inverter  inverter_0
timestamp 1700276902
transform 1 0 50980 0 1 145
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1700276902
transform 1 0 7480 0 1 145
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1700276902
transform 1 0 14730 0 1 145
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1700276902
transform 1 0 21980 0 1 145
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1700276902
transform 1 0 29230 0 1 145
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1700276902
transform 1 0 36480 0 1 145
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1700276902
transform 1 0 43730 0 1 145
box -240 -145 -30 185
use ladder  ladder_0
timestamp 1700206437
transform 1 0 10310 0 1 985
box -10460 -640 48210 205
<< end >>
