magic
tech sky130A
timestamp 1700276151
<< nwell >>
rect -3520 -105 18450 1530
<< nmos >>
rect 19700 -50 20500 1150
rect 21300 -50 22100 1150
rect 22900 -50 23700 1150
rect 24500 -50 25300 1150
rect 26100 -50 26900 1150
rect -2320 -1545 -1520 -345
rect -720 -1545 80 -345
rect 1801 -1545 2601 -345
rect 3401 -1545 4201 -345
rect 5001 -1545 5801 -345
rect 6601 -1545 7401 -345
rect 8201 -1545 9001 -345
rect 9801 -1545 10601 -345
rect 11401 -1545 12201 -345
rect 13001 -1545 13801 -345
rect 14601 -1545 15401 -345
rect 16201 -1545 17001 -345
rect 17801 -1545 18601 -345
rect 19401 -1545 20201 -345
rect 21001 -1545 21801 -345
rect 22601 -1545 23401 -345
rect 24201 -1545 25001 -345
rect 25801 -1545 26601 -345
rect 28296 -1545 29096 -345
rect 29896 -1545 30696 -345
<< pmos >>
rect -2315 -50 -1515 1150
rect -715 -50 85 1150
rect 885 -50 1685 1150
rect 2485 -50 3285 1150
rect 4085 -50 4885 1150
rect 6645 -50 7445 1150
rect 8245 -50 9045 1150
rect 10800 -50 11600 1150
rect 12400 -50 13200 1150
rect 15050 -50 15850 1150
rect 16650 -50 17450 1150
<< ndiff >>
rect 18900 1050 19700 1150
rect 18900 50 19000 1050
rect 19600 50 19700 1050
rect 18900 -50 19700 50
rect 20500 1050 21300 1150
rect 20500 50 20600 1050
rect 21200 50 21300 1050
rect 20500 -50 21300 50
rect 22100 1050 22900 1150
rect 22100 50 22200 1050
rect 22800 50 22900 1050
rect 22100 -50 22900 50
rect 23700 1050 24500 1150
rect 23700 50 23800 1050
rect 24400 50 24500 1050
rect 23700 -50 24500 50
rect 25300 1050 26100 1150
rect 25300 50 25400 1050
rect 26000 50 26100 1050
rect 25300 -50 26100 50
rect 26900 1100 27700 1150
rect 26900 1050 27650 1100
rect 26900 50 27000 1050
rect 27600 50 27650 1050
rect 26900 0 27650 50
rect 26900 -50 27700 0
rect -3120 -445 -2320 -345
rect -3120 -1445 -3020 -445
rect -2420 -1445 -2320 -445
rect -3120 -1545 -2320 -1445
rect -1520 -445 -720 -345
rect -1520 -1445 -1420 -445
rect -820 -1445 -720 -445
rect -1520 -1545 -720 -1445
rect 80 -445 880 -345
rect 80 -1445 180 -445
rect 780 -1445 880 -445
rect 80 -1545 880 -1445
rect 1001 -445 1801 -345
rect 1001 -1445 1101 -445
rect 1701 -1445 1801 -445
rect 1001 -1545 1801 -1445
rect 2601 -445 3401 -345
rect 2601 -1445 2701 -445
rect 3301 -1445 3401 -445
rect 2601 -1545 3401 -1445
rect 4201 -445 5001 -345
rect 4201 -1445 4301 -445
rect 4901 -1445 5001 -445
rect 4201 -1545 5001 -1445
rect 5801 -445 6601 -345
rect 5801 -1445 5901 -445
rect 6501 -1445 6601 -445
rect 5801 -1545 6601 -1445
rect 7401 -445 8201 -345
rect 7401 -1445 7501 -445
rect 8101 -1445 8201 -445
rect 7401 -1545 8201 -1445
rect 9001 -445 9801 -345
rect 9001 -1445 9101 -445
rect 9701 -1445 9801 -445
rect 9001 -1545 9801 -1445
rect 10601 -445 11401 -345
rect 10601 -1445 10701 -445
rect 11301 -1445 11401 -445
rect 10601 -1545 11401 -1445
rect 12201 -445 13001 -345
rect 12201 -1445 12301 -445
rect 12901 -1445 13001 -445
rect 12201 -1545 13001 -1445
rect 13801 -445 14601 -345
rect 13801 -1445 13901 -445
rect 14501 -1445 14601 -445
rect 13801 -1545 14601 -1445
rect 15401 -445 16201 -345
rect 15401 -1445 15501 -445
rect 16101 -1445 16201 -445
rect 15401 -1545 16201 -1445
rect 17001 -445 17801 -345
rect 17001 -1445 17101 -445
rect 17701 -1445 17801 -445
rect 17001 -1545 17801 -1445
rect 18601 -445 19401 -345
rect 18601 -1445 18701 -445
rect 19301 -1445 19401 -445
rect 18601 -1545 19401 -1445
rect 20201 -445 21001 -345
rect 20201 -1445 20301 -445
rect 20901 -1445 21001 -445
rect 20201 -1545 21001 -1445
rect 21801 -445 22601 -345
rect 21801 -1445 21901 -445
rect 22501 -1445 22601 -445
rect 21801 -1545 22601 -1445
rect 23401 -445 24201 -345
rect 23401 -1445 23501 -445
rect 24101 -1445 24201 -445
rect 23401 -1545 24201 -1445
rect 25001 -445 25801 -345
rect 25001 -1445 25101 -445
rect 25701 -1445 25801 -445
rect 25001 -1545 25801 -1445
rect 26601 -445 27400 -345
rect 26601 -1445 26701 -445
rect 27301 -1445 27400 -445
rect 26601 -1545 27400 -1445
rect 27496 -445 28296 -345
rect 27496 -1445 27596 -445
rect 28196 -1445 28296 -445
rect 27496 -1545 28296 -1445
rect 29096 -445 29896 -345
rect 29096 -1445 29195 -445
rect 29795 -1445 29896 -445
rect 29096 -1545 29896 -1445
rect 30696 -445 31495 -345
rect 30696 -1445 30796 -445
rect 31396 -1445 31495 -445
rect 30696 -1545 31495 -1445
<< pdiff >>
rect -3115 1050 -2315 1150
rect -3115 50 -3015 1050
rect -2415 50 -2315 1050
rect -3115 -50 -2315 50
rect -1515 1050 -715 1150
rect -1515 50 -1415 1050
rect -815 50 -715 1050
rect -1515 -50 -715 50
rect 85 1050 885 1150
rect 85 50 185 1050
rect 785 50 885 1050
rect 85 -50 885 50
rect 1685 1050 2485 1150
rect 1685 50 1785 1050
rect 2385 50 2485 1050
rect 1685 -50 2485 50
rect 3285 1050 4085 1150
rect 3285 50 3385 1050
rect 3985 50 4085 1050
rect 3285 -50 4085 50
rect 4885 1050 5685 1150
rect 4885 50 4985 1050
rect 5585 50 5685 1050
rect 4885 -50 5685 50
rect 5845 1050 6645 1150
rect 5845 50 5945 1050
rect 6545 50 6645 1050
rect 5845 -50 6645 50
rect 7445 1050 8245 1150
rect 7445 50 7545 1050
rect 8145 50 8245 1050
rect 7445 -50 8245 50
rect 9045 1050 9845 1150
rect 9045 50 9145 1050
rect 9745 50 9845 1050
rect 9045 -50 9845 50
rect 10000 1050 10800 1150
rect 10000 50 10100 1050
rect 10700 50 10800 1050
rect 10000 -50 10800 50
rect 11600 1050 12400 1150
rect 11600 50 11700 1050
rect 12300 50 12400 1050
rect 11600 -50 12400 50
rect 13200 1050 14000 1150
rect 13200 50 13300 1050
rect 13900 50 14000 1050
rect 13200 -50 14000 50
rect 14250 1050 15050 1150
rect 14250 50 14350 1050
rect 14950 50 15050 1050
rect 14250 -50 15050 50
rect 15850 1050 16650 1150
rect 15850 50 15950 1050
rect 16550 50 16650 1050
rect 15850 -50 16650 50
rect 17450 1050 18250 1150
rect 17450 50 17550 1050
rect 18150 50 18250 1050
rect 17450 -50 18250 50
<< ndiffc >>
rect 19000 50 19600 1050
rect 20600 50 21200 1050
rect 22200 50 22800 1050
rect 23800 50 24400 1050
rect 25400 50 26000 1050
rect 27000 50 27600 1050
rect -3020 -1445 -2420 -445
rect -1420 -1445 -820 -445
rect 180 -1445 780 -445
rect 1101 -1445 1701 -445
rect 2701 -1445 3301 -445
rect 4301 -1445 4901 -445
rect 5901 -1445 6501 -445
rect 7501 -1445 8101 -445
rect 9101 -1445 9701 -445
rect 10701 -1445 11301 -445
rect 12301 -1445 12901 -445
rect 13901 -1445 14501 -445
rect 15501 -1445 16101 -445
rect 17101 -1445 17701 -445
rect 18701 -1445 19301 -445
rect 20301 -1445 20901 -445
rect 21901 -1445 22501 -445
rect 23501 -1445 24101 -445
rect 25101 -1445 25701 -445
rect 26701 -1445 27301 -445
rect 27596 -1445 28196 -445
rect 29195 -1445 29795 -445
rect 30796 -1445 31396 -445
<< pdiffc >>
rect -3015 50 -2415 1050
rect -1415 50 -815 1050
rect 185 50 785 1050
rect 1785 50 2385 1050
rect 3385 50 3985 1050
rect 4985 50 5585 1050
rect 5945 50 6545 1050
rect 7545 50 8145 1050
rect 9145 50 9745 1050
rect 10100 50 10700 1050
rect 11700 50 12300 1050
rect 13300 50 13900 1050
rect 14350 50 14950 1050
rect 15950 50 16550 1050
rect 17550 50 18150 1050
<< psubdiff >>
rect 20300 1350 20600 1400
rect 20300 1300 20350 1350
rect 20550 1300 20600 1350
rect 20300 1250 20600 1300
rect 23350 1350 23650 1400
rect 23350 1300 23400 1350
rect 23600 1300 23650 1350
rect 23350 1250 23650 1300
rect 25850 1350 26150 1400
rect 25850 1300 25900 1350
rect 26100 1300 26150 1350
rect 25850 1250 26150 1300
rect 27700 1100 28000 1150
rect 27650 1050 28000 1100
rect 27650 50 27750 1050
rect 27900 50 28000 1050
rect 27650 0 28000 50
rect 27700 -50 28000 0
rect -3420 -445 -3120 -345
rect -3420 -1445 -3320 -445
rect -3170 -1445 -3120 -445
rect -3420 -1545 -3120 -1445
rect 31495 -445 31795 -345
rect 31495 -1445 31545 -445
rect 31695 -1445 31795 -445
rect 31495 -1545 31795 -1445
rect -1220 -1660 -920 -1610
rect -1220 -1710 -1170 -1660
rect -970 -1710 -920 -1660
rect -1220 -1760 -920 -1710
rect 1101 -1660 1401 -1610
rect 1101 -1710 1151 -1660
rect 1351 -1710 1401 -1660
rect 1101 -1760 1401 -1710
rect 4101 -1660 4401 -1610
rect 4101 -1710 4151 -1660
rect 4351 -1710 4401 -1660
rect 4101 -1760 4401 -1710
rect 7101 -1660 7401 -1610
rect 7101 -1710 7151 -1660
rect 7351 -1710 7401 -1660
rect 7101 -1760 7401 -1710
rect 10101 -1660 10401 -1610
rect 10101 -1710 10151 -1660
rect 10351 -1710 10401 -1660
rect 10101 -1760 10401 -1710
rect 13101 -1660 13401 -1610
rect 13101 -1710 13151 -1660
rect 13351 -1710 13401 -1660
rect 13101 -1760 13401 -1710
rect 16101 -1660 16401 -1610
rect 16101 -1710 16151 -1660
rect 16351 -1710 16401 -1660
rect 16101 -1760 16401 -1710
rect 19601 -1660 19901 -1610
rect 19601 -1710 19651 -1660
rect 19851 -1710 19901 -1660
rect 19601 -1760 19901 -1710
rect 22601 -1660 22901 -1610
rect 22601 -1710 22651 -1660
rect 22851 -1710 22901 -1660
rect 22601 -1760 22901 -1710
rect 25801 -1660 26101 -1610
rect 25801 -1710 25851 -1660
rect 26051 -1710 26101 -1660
rect 25801 -1760 26101 -1710
rect 28161 -1660 28461 -1610
rect 28161 -1710 28211 -1660
rect 28411 -1710 28461 -1660
rect 28161 -1760 28461 -1710
<< nsubdiff >>
rect -1395 1350 -1095 1400
rect -1395 1300 -1345 1350
rect -1145 1300 -1095 1350
rect -1395 1250 -1095 1300
rect 1785 1350 2085 1400
rect 1785 1300 1835 1350
rect 2035 1300 2085 1350
rect 1785 1250 2085 1300
rect 4785 1350 5085 1400
rect 4785 1300 4835 1350
rect 5035 1300 5085 1350
rect 4785 1250 5085 1300
rect 7695 1350 7995 1400
rect 7695 1300 7745 1350
rect 7945 1300 7995 1350
rect 7695 1250 7995 1300
rect 10600 1350 10900 1400
rect 10600 1300 10650 1350
rect 10850 1300 10900 1350
rect 10600 1250 10900 1300
rect 13600 1350 13900 1400
rect 13600 1300 13650 1350
rect 13850 1300 13900 1350
rect 13600 1250 13900 1300
rect 16600 1350 16900 1400
rect 16600 1300 16650 1350
rect 16850 1300 16900 1350
rect 16600 1250 16900 1300
rect -3415 1050 -3115 1150
rect -3415 50 -3315 1050
rect -3165 50 -3115 1050
rect -3415 -50 -3115 50
<< psubdiffcont >>
rect 20350 1300 20550 1350
rect 23400 1300 23600 1350
rect 25900 1300 26100 1350
rect 27750 50 27900 1050
rect -3320 -1445 -3170 -445
rect 31545 -1445 31695 -445
rect -1170 -1710 -970 -1660
rect 1151 -1710 1351 -1660
rect 4151 -1710 4351 -1660
rect 7151 -1710 7351 -1660
rect 10151 -1710 10351 -1660
rect 13151 -1710 13351 -1660
rect 16151 -1710 16351 -1660
rect 19651 -1710 19851 -1660
rect 22651 -1710 22851 -1660
rect 25851 -1710 26051 -1660
rect 28211 -1710 28411 -1660
<< nsubdiffcont >>
rect -1345 1300 -1145 1350
rect 1835 1300 2035 1350
rect 4835 1300 5035 1350
rect 7745 1300 7945 1350
rect 10650 1300 10850 1350
rect 13650 1300 13850 1350
rect 16650 1300 16850 1350
rect -3315 50 -3165 1050
<< poly >>
rect -2315 1250 -1515 1265
rect 6645 1250 7445 1265
rect -2315 1195 -2300 1250
rect -1530 1195 -1515 1250
rect -2315 1150 -1515 1195
rect -715 1150 85 1200
rect 885 1150 1685 1200
rect 2485 1150 3285 1205
rect 4085 1150 4885 1200
rect 6645 1195 6660 1250
rect 7435 1195 7445 1250
rect 6645 1150 7445 1195
rect 8245 1150 9045 1200
rect 10800 1150 11600 1200
rect 12400 1150 13200 1200
rect 15050 1150 15850 1200
rect 16650 1150 17450 1200
rect 19700 1150 20500 1200
rect 21300 1150 22100 1200
rect 22900 1150 23700 1200
rect 24500 1150 25300 1200
rect 26100 1150 26900 1200
rect -2315 -100 -1515 -50
rect -715 -100 85 -50
rect 885 -100 1685 -50
rect 2485 -100 3285 -50
rect 4085 -100 4885 -50
rect -715 -115 4885 -100
rect -715 -150 2495 -115
rect 2480 -170 2495 -150
rect 3270 -150 4885 -115
rect 6645 -100 7445 -50
rect 8245 -100 9045 -50
rect 10800 -100 11600 -50
rect 12400 -100 13200 -50
rect 15050 -100 15850 -50
rect 16650 -100 17450 -50
rect 6645 -105 17450 -100
rect 18740 -80 19540 -65
rect 18740 -105 18755 -80
rect 6645 -135 18755 -105
rect 19525 -135 19540 -80
rect 6645 -150 19540 -135
rect 19700 -100 20500 -50
rect 21300 -100 22100 -50
rect 22900 -100 23700 -50
rect 24500 -100 25300 -50
rect 19700 -115 25300 -100
rect 19700 -150 21315 -115
rect 3270 -170 3285 -150
rect 2480 -185 3285 -170
rect 21300 -170 21315 -150
rect 22085 -150 25300 -115
rect 26100 -115 26900 -50
rect 22085 -170 22100 -150
rect 21300 -185 22100 -170
rect 26100 -170 26115 -115
rect 26885 -170 26900 -115
rect 26100 -185 26900 -170
rect 11400 -220 12200 -205
rect 11400 -245 11415 -220
rect -720 -275 11415 -245
rect 12185 -245 12200 -220
rect 12185 -275 29095 -245
rect -720 -295 29095 -275
rect -2320 -345 -1520 -295
rect -720 -345 80 -295
rect 1801 -345 2601 -295
rect 3401 -345 4201 -295
rect 5001 -345 5801 -295
rect 6601 -345 7401 -295
rect 8201 -345 9001 -295
rect 9801 -345 10601 -295
rect 11401 -345 12201 -295
rect 13001 -345 13801 -295
rect 14601 -345 15401 -295
rect 16201 -345 17001 -295
rect 17801 -345 18601 -295
rect 19401 -345 20201 -295
rect 21001 -345 21801 -295
rect 22601 -345 23401 -295
rect 24201 -345 25001 -295
rect 25801 -345 26601 -295
rect 28296 -345 29096 -295
rect 29896 -345 30696 -295
rect -2320 -1600 -1520 -1545
rect -720 -1595 80 -1545
rect 1801 -1595 2601 -1545
rect 3401 -1595 4201 -1545
rect 5001 -1595 5801 -1545
rect 6601 -1595 7401 -1545
rect 8201 -1595 9001 -1545
rect 9801 -1595 10601 -1545
rect 11401 -1595 12201 -1545
rect 13001 -1595 13801 -1545
rect 14601 -1595 15401 -1545
rect 16201 -1595 17001 -1545
rect 17801 -1595 18601 -1545
rect 19401 -1595 20201 -1545
rect 21001 -1595 21801 -1545
rect 22601 -1595 23401 -1545
rect 24201 -1595 25001 -1545
rect 25801 -1595 26601 -1545
rect 28296 -1595 29096 -1545
rect 29896 -1595 30696 -1545
rect -2320 -1655 -2305 -1600
rect -1535 -1655 -1520 -1600
rect -2320 -1670 -1520 -1655
rect 900 -1630 1045 -1605
rect 29895 -1610 30695 -1595
rect 900 -1720 925 -1630
rect 1020 -1720 1045 -1630
rect 900 -1745 1045 -1720
rect 900 -1785 940 -1745
rect 29895 -1665 29910 -1610
rect 30680 -1665 30695 -1610
rect 29895 -1680 30695 -1665
rect -3520 -1825 940 -1785
<< polycont >>
rect -2300 1195 -1530 1250
rect 6660 1195 7435 1250
rect 2495 -170 3270 -115
rect 18755 -135 19525 -80
rect 21315 -170 22085 -115
rect 26115 -170 26885 -115
rect 11415 -275 12185 -220
rect -2305 -1655 -1535 -1600
rect 925 -1720 1020 -1630
rect 29910 -1665 30680 -1610
<< locali >>
rect -3520 1435 9795 1485
rect -1370 1350 -1115 1375
rect -1370 1300 -1345 1350
rect -1145 1300 -1115 1350
rect -1370 1280 -1115 1300
rect 1810 1350 2065 1375
rect 1810 1300 1835 1350
rect 2035 1300 2065 1350
rect 1810 1280 2065 1300
rect 4810 1350 5065 1375
rect 4810 1300 4835 1350
rect 5035 1300 5065 1350
rect 4810 1280 5065 1300
rect 7720 1350 7975 1375
rect 7720 1300 7745 1350
rect 7945 1300 7975 1350
rect 7720 1280 7975 1300
rect -2315 1250 -1515 1265
rect -2315 1195 -2300 1250
rect -1530 1195 -1515 1250
rect 6645 1250 7445 1265
rect 6645 1215 6660 1250
rect -2315 1180 -1515 1195
rect -1465 1195 6660 1215
rect 7435 1195 7445 1250
rect -1465 1180 7445 1195
rect -3365 1050 -2365 1100
rect -3365 50 -3315 1050
rect -3165 50 -3015 1050
rect -2415 50 -2365 1050
rect -3365 0 -2365 50
rect -1465 1050 -765 1180
rect -1465 50 -1415 1050
rect -815 50 -765 1050
rect -1465 -85 -765 50
rect 135 1050 835 1100
rect 135 50 185 1050
rect 785 50 835 1050
rect 135 0 835 50
rect 1735 1050 2435 1105
rect 1735 50 1785 1050
rect 2385 50 2435 1050
rect -3520 -130 -765 -85
rect 1735 -100 2435 50
rect 3335 1050 4035 1100
rect 3335 50 3385 1050
rect 3985 50 4035 1050
rect 3335 0 4035 50
rect 4935 1050 5635 1180
rect 4935 50 4985 1050
rect 5585 50 5635 1050
rect 4935 0 5635 50
rect 5895 1050 6595 1100
rect 5895 50 5945 1050
rect 6545 50 6595 1050
rect 5895 0 6595 50
rect 7495 1050 8195 1100
rect 7495 50 7545 1050
rect 8145 50 8195 1050
rect 7495 0 8195 50
rect 9095 1050 9795 1435
rect 10625 1350 10880 1375
rect 10625 1300 10650 1350
rect 10850 1300 10880 1350
rect 10625 1280 10880 1300
rect 13625 1350 13880 1375
rect 13625 1300 13650 1350
rect 13850 1300 13880 1350
rect 13625 1280 13880 1300
rect 16625 1350 16880 1375
rect 16625 1300 16650 1350
rect 16850 1300 16880 1350
rect 16625 1280 16880 1300
rect 20325 1350 20580 1375
rect 20325 1300 20350 1350
rect 20550 1300 20580 1350
rect 20325 1280 20580 1300
rect 23375 1350 23630 1375
rect 23375 1300 23400 1350
rect 23600 1300 23630 1350
rect 23375 1280 23630 1300
rect 25875 1350 26130 1375
rect 25875 1300 25900 1350
rect 26100 1300 26130 1350
rect 25875 1280 26130 1300
rect 22150 1210 22850 1215
rect 11650 1160 22850 1210
rect 9095 50 9145 1050
rect 9745 50 9795 1050
rect 1735 -115 3285 -100
rect 1735 -150 2495 -115
rect 1735 -210 2435 -150
rect 2480 -170 2495 -150
rect 3270 -170 3285 -115
rect 2480 -185 3285 -170
rect 5945 -185 6590 0
rect 9095 -45 9795 50
rect 10050 1050 10750 1100
rect 10050 50 10100 1050
rect 10700 50 10750 1050
rect 10050 0 10750 50
rect 11650 1050 12350 1160
rect 11650 50 11700 1050
rect 12300 50 12350 1050
rect 11650 0 12350 50
rect 13250 1050 13950 1100
rect 13250 50 13300 1050
rect 13900 50 13950 1050
rect 13250 0 13950 50
rect 14300 1050 15000 1100
rect 14300 50 14350 1050
rect 14950 50 15000 1050
rect 14300 0 15000 50
rect 15900 1050 16600 1100
rect 15900 50 15950 1050
rect 16550 50 16600 1050
rect 15900 0 16600 50
rect 17500 1050 18200 1100
rect 17500 50 17550 1050
rect 18150 50 18200 1050
rect 9095 -75 9800 -45
rect 9100 -85 9800 -75
rect 14305 -85 14995 0
rect 9100 -130 14995 -85
rect 17500 -185 18200 50
rect 18950 1050 19650 1100
rect 18950 50 19000 1050
rect 19600 50 19650 1050
rect 18950 0 19650 50
rect 20550 1050 21250 1100
rect 20550 50 20600 1050
rect 21200 50 21250 1050
rect 20550 0 21250 50
rect 22150 1050 22850 1160
rect 22150 50 22200 1050
rect 22800 50 22850 1050
rect 18950 -65 19540 0
rect 18740 -80 19540 -65
rect 18740 -135 18755 -80
rect 19525 -135 19540 -80
rect 22150 -100 22850 50
rect 23750 1050 24450 1100
rect 23750 50 23800 1050
rect 24400 50 24450 1050
rect 23750 0 24450 50
rect 25350 1050 26050 1100
rect 25350 50 25400 1050
rect 26000 50 26050 1050
rect 25350 0 26050 50
rect 26950 1050 27950 1100
rect 26950 50 27000 1050
rect 27600 50 27750 1050
rect 27900 50 27950 1050
rect 26950 0 27950 50
rect 18740 -150 19540 -135
rect 1550 -265 2250 -210
rect 5945 -220 18200 -185
rect 5945 -235 11415 -220
rect -1470 -310 2250 -265
rect 11400 -275 11415 -235
rect 12185 -235 18200 -220
rect 19495 -210 19540 -150
rect 21300 -115 22855 -100
rect 21300 -170 21315 -115
rect 22085 -150 22855 -115
rect 22085 -170 22100 -150
rect 21300 -185 22100 -170
rect 25350 -210 26005 0
rect 26100 -115 26900 -100
rect 26100 -170 26115 -115
rect 26885 -170 26900 -115
rect 26100 -185 26900 -170
rect 12185 -275 12200 -235
rect 19495 -240 26005 -210
rect 11400 -295 12200 -275
rect -1470 -395 -765 -310
rect 2650 -345 25745 -295
rect 2650 -395 3350 -345
rect 5850 -395 6555 -345
rect 9050 -395 9750 -345
rect 12250 -395 12950 -345
rect 15450 -395 16150 -345
rect 18650 -395 19350 -345
rect 21850 -395 22550 -345
rect 25050 -395 25745 -345
rect -3370 -445 -2370 -395
rect -3370 -1445 -3320 -445
rect -3170 -1445 -3020 -445
rect -2420 -1445 -2370 -445
rect -3370 -1495 -2370 -1445
rect -1470 -445 -770 -395
rect -1470 -1445 -1420 -445
rect -820 -1445 -770 -445
rect -1470 -1495 -770 -1445
rect 130 -445 830 -395
rect 130 -1445 180 -445
rect 780 -1445 830 -445
rect 130 -1495 830 -1445
rect 1051 -445 1751 -395
rect 1051 -1445 1101 -445
rect 1701 -1445 1751 -445
rect 1051 -1495 1751 -1445
rect 2651 -445 3351 -395
rect 2651 -1445 2701 -445
rect 3301 -1445 3351 -445
rect 2651 -1495 3351 -1445
rect 4251 -445 4951 -395
rect 4251 -1445 4301 -445
rect 4901 -1445 4951 -445
rect 4251 -1495 4951 -1445
rect 5851 -445 6551 -395
rect 5851 -1445 5901 -445
rect 6501 -1445 6551 -445
rect 5851 -1495 6551 -1445
rect 7451 -445 8151 -395
rect 7451 -1445 7501 -445
rect 8101 -1445 8151 -445
rect 7451 -1495 8151 -1445
rect 9051 -445 9751 -395
rect 9051 -1445 9101 -445
rect 9701 -1445 9751 -445
rect 9051 -1495 9751 -1445
rect 10651 -445 11351 -395
rect 12250 -400 12951 -395
rect 10651 -1445 10701 -445
rect 11301 -1445 11351 -445
rect 10651 -1495 11351 -1445
rect 12251 -445 12951 -400
rect 12251 -1445 12301 -445
rect 12901 -1445 12951 -445
rect 12251 -1495 12951 -1445
rect 13851 -445 14551 -395
rect 13851 -1445 13901 -445
rect 14501 -1445 14551 -445
rect 13851 -1495 14551 -1445
rect 15451 -445 16151 -395
rect 15451 -1445 15501 -445
rect 16101 -1445 16151 -445
rect 15451 -1495 16151 -1445
rect 17051 -445 17751 -395
rect 17051 -1445 17101 -445
rect 17701 -1445 17751 -445
rect 17051 -1495 17751 -1445
rect 18651 -445 19351 -395
rect 18651 -1445 18701 -445
rect 19301 -1445 19351 -445
rect 18651 -1495 19351 -1445
rect 20251 -445 20951 -395
rect 20251 -1445 20301 -445
rect 20901 -1445 20951 -445
rect 20251 -1495 20951 -1445
rect 21851 -445 22551 -395
rect 21851 -1445 21901 -445
rect 22501 -1445 22551 -445
rect 21851 -1495 22551 -1445
rect 23451 -445 24151 -395
rect 23451 -1445 23501 -445
rect 24101 -1445 24151 -445
rect 23451 -1495 24151 -1445
rect 25051 -445 25751 -395
rect 25051 -1445 25101 -445
rect 25701 -1445 25751 -445
rect 25051 -1495 25751 -1445
rect 26651 -410 27350 -395
rect 26651 -445 27351 -410
rect 26651 -1445 26701 -445
rect 27301 -1445 27351 -445
rect 26651 -1495 27351 -1445
rect 27496 -445 28246 -395
rect 27496 -1445 27596 -445
rect 28196 -1445 28246 -445
rect 29146 -445 29846 -395
rect 29146 -1440 29195 -445
rect 27496 -1495 28246 -1445
rect 29145 -1445 29195 -1440
rect 29795 -1445 29846 -445
rect 29145 -1495 29846 -1445
rect 30746 -445 31745 -395
rect 30746 -1445 30796 -445
rect 31396 -1445 31545 -445
rect 31695 -1445 31745 -445
rect 30746 -1495 31745 -1445
rect -2320 -1600 -1520 -1585
rect -2320 -1655 -2305 -1600
rect -1535 -1655 -1520 -1600
rect -2320 -1670 -1520 -1655
rect -1470 -1775 -1420 -1495
rect 1050 -1535 1750 -1495
rect 4250 -1535 4950 -1495
rect 7450 -1535 8150 -1495
rect 10650 -1535 11350 -1495
rect 13850 -1535 14550 -1495
rect 17050 -1535 17750 -1495
rect 20250 -1535 20950 -1495
rect 23450 -1535 24150 -1495
rect 26650 -1535 27350 -1495
rect 1000 -1585 27350 -1535
rect 1000 -1605 1045 -1585
rect 29145 -1590 29845 -1495
rect 31445 -1496 31490 -1495
rect 900 -1630 1045 -1605
rect -1195 -1660 -940 -1635
rect -1195 -1710 -1170 -1660
rect -970 -1710 -940 -1660
rect -1195 -1730 -940 -1710
rect 900 -1720 925 -1630
rect 1020 -1720 1045 -1630
rect 900 -1745 1045 -1720
rect 1126 -1660 1381 -1635
rect 1126 -1710 1151 -1660
rect 1351 -1710 1381 -1660
rect 1126 -1730 1381 -1710
rect 4126 -1660 4381 -1635
rect 4126 -1710 4151 -1660
rect 4351 -1710 4381 -1660
rect 4126 -1730 4381 -1710
rect 7126 -1660 7381 -1635
rect 7126 -1710 7151 -1660
rect 7351 -1710 7381 -1660
rect 7126 -1730 7381 -1710
rect 10126 -1660 10381 -1635
rect 10126 -1710 10151 -1660
rect 10351 -1710 10381 -1660
rect 10126 -1730 10381 -1710
rect 13126 -1660 13381 -1635
rect 13126 -1710 13151 -1660
rect 13351 -1710 13381 -1660
rect 13126 -1730 13381 -1710
rect 16126 -1660 16381 -1635
rect 16126 -1710 16151 -1660
rect 16351 -1710 16381 -1660
rect 16126 -1730 16381 -1710
rect 19626 -1660 19881 -1635
rect 19626 -1710 19651 -1660
rect 19851 -1710 19881 -1660
rect 19626 -1730 19881 -1710
rect 22626 -1660 22881 -1635
rect 22626 -1710 22651 -1660
rect 22851 -1710 22881 -1660
rect 22626 -1730 22881 -1710
rect 25826 -1660 26081 -1635
rect 25826 -1710 25851 -1660
rect 26051 -1710 26081 -1660
rect 25826 -1730 26081 -1710
rect 28186 -1660 28441 -1635
rect 28186 -1710 28211 -1660
rect 28411 -1710 28441 -1660
rect 28186 -1730 28441 -1710
rect 29745 -1775 29795 -1590
rect 29895 -1610 30695 -1595
rect 29895 -1665 29910 -1610
rect 30680 -1665 30695 -1610
rect 29895 -1680 30695 -1665
rect -1470 -1825 29795 -1775
<< viali >>
rect -1345 1300 -1145 1350
rect 1835 1300 2035 1350
rect 4835 1300 5035 1350
rect 7745 1300 7945 1350
rect -2300 1195 -1530 1250
rect -3315 50 -3165 1050
rect -3015 50 -2415 1050
rect 185 50 785 1050
rect 3385 50 3985 1050
rect 7545 50 8145 1050
rect 10650 1300 10850 1350
rect 13650 1300 13850 1350
rect 16650 1300 16850 1350
rect 20350 1300 20550 1350
rect 23400 1300 23600 1350
rect 25900 1300 26100 1350
rect 10100 50 10700 1050
rect 13300 50 13900 1050
rect 15950 50 16550 1050
rect 20600 50 21200 1050
rect 23800 50 24400 1050
rect 27000 50 27600 1050
rect 27750 50 27900 1050
rect 26115 -170 26885 -115
rect -3320 -1445 -3170 -445
rect -3020 -1445 -2420 -445
rect 180 -1445 780 -445
rect 27596 -1445 28196 -445
rect 30796 -1445 31396 -445
rect 31545 -1445 31695 -445
rect -2305 -1655 -1535 -1600
rect -1170 -1710 -970 -1660
rect 1151 -1710 1351 -1660
rect 4151 -1710 4351 -1660
rect 7151 -1710 7351 -1660
rect 10151 -1710 10351 -1660
rect 13151 -1710 13351 -1660
rect 16151 -1710 16351 -1660
rect 19651 -1710 19851 -1660
rect 22651 -1710 22851 -1660
rect 25851 -1710 26051 -1660
rect 28211 -1710 28411 -1660
rect 29910 -1665 30680 -1610
<< metal1 >>
rect -3520 1350 18450 1450
rect -3520 1300 -1345 1350
rect -1145 1300 1835 1350
rect 2035 1300 4835 1350
rect 5035 1300 7745 1350
rect 7945 1300 10650 1350
rect 10850 1300 13650 1350
rect 13850 1300 16650 1350
rect 16850 1300 18450 1350
rect -3520 1250 18450 1300
rect -3520 1195 -2300 1250
rect -1530 1195 18450 1250
rect -3520 1050 18450 1195
rect -3520 50 -3315 1050
rect -3165 50 -3015 1050
rect -2415 50 185 1050
rect 785 50 3385 1050
rect 3985 50 7545 1050
rect 8145 50 10100 1050
rect 10700 50 13300 1050
rect 13900 50 15950 1050
rect 16550 50 18450 1050
rect -3520 -15 18450 50
rect 18900 1350 28100 1450
rect 18900 1300 20350 1350
rect 20550 1300 23400 1350
rect 23600 1300 25900 1350
rect 26100 1300 28100 1350
rect 18900 1050 28100 1300
rect 18900 50 20600 1050
rect 21200 50 23800 1050
rect 24400 50 27000 1050
rect 27600 50 27750 1050
rect 27900 50 28100 1050
rect 18900 -115 28100 50
rect 18900 -170 26115 -115
rect 26885 -170 28100 -115
rect 18900 -395 28100 -170
rect -3520 -445 31825 -395
rect -3520 -1445 -3320 -445
rect -3170 -1445 -3020 -445
rect -2420 -1445 180 -445
rect 780 -1445 27596 -445
rect 28196 -1445 30796 -445
rect 31396 -1445 31545 -445
rect 31695 -1445 31825 -445
rect -3520 -1600 31825 -1445
rect -3520 -1655 -2305 -1600
rect -1535 -1610 31825 -1600
rect -1535 -1655 29910 -1610
rect -3520 -1660 29910 -1655
rect -3520 -1710 -1170 -1660
rect -970 -1710 1151 -1660
rect 1351 -1710 4151 -1660
rect 4351 -1710 7151 -1660
rect 7351 -1710 10151 -1660
rect 10351 -1710 13151 -1660
rect 13351 -1710 16151 -1660
rect 16351 -1710 19651 -1660
rect 19851 -1710 22651 -1660
rect 22851 -1710 25851 -1660
rect 26051 -1710 28211 -1660
rect 28411 -1665 29910 -1660
rect 30680 -1665 31825 -1610
rect 28411 -1710 31825 -1665
rect -3520 -1760 31825 -1710
<< labels >>
rlabel locali -3520 1460 -3520 1460 7 Iin
port 1 w
rlabel locali -3520 -110 -3520 -110 7 Vbp
port 2 w
rlabel poly -3520 -1805 -3520 -1805 7 Ires
port 3 w
rlabel metal1 -3520 545 -3520 545 7 VP
port 4 w
rlabel metal1 -3520 -945 -3520 -945 7 VN
port 5 w
<< end >>
