magic
tech sky130A
timestamp 1700269757
<< psubdiff >>
rect 3200 1285 3300 1300
rect 3200 1265 3215 1285
rect 3285 1265 3300 1285
rect 3200 1250 3300 1265
rect 5200 1285 5300 1300
rect 5200 1265 5215 1285
rect 5285 1265 5300 1285
rect 5200 1250 5300 1265
rect 7200 1285 7300 1300
rect 7200 1265 7215 1285
rect 7285 1265 7300 1285
rect 7200 1250 7300 1265
rect 9200 1285 9300 1300
rect 9200 1265 9215 1285
rect 9285 1265 9300 1285
rect 9200 1250 9300 1265
rect 11200 1285 11300 1300
rect 11200 1265 11215 1285
rect 11285 1265 11300 1285
rect 11200 1250 11300 1265
rect 13200 1285 13300 1300
rect 13200 1265 13215 1285
rect 13285 1265 13300 1285
rect 13200 1250 13300 1265
rect 15200 1285 15300 1300
rect 15200 1265 15215 1285
rect 15285 1265 15300 1285
rect 15200 1250 15300 1265
rect 17200 1285 17300 1300
rect 17200 1265 17215 1285
rect 17285 1265 17300 1285
rect 17200 1250 17300 1265
rect 19200 1285 19300 1300
rect 19200 1265 19215 1285
rect 19285 1265 19300 1285
rect 19200 1250 19300 1265
rect 21200 1285 21300 1300
rect 21200 1265 21215 1285
rect 21285 1265 21300 1285
rect 21200 1250 21300 1265
rect 23200 1285 23300 1300
rect 23200 1265 23215 1285
rect 23285 1265 23300 1285
rect 23200 1250 23300 1265
rect 25200 1285 25300 1300
rect 25200 1265 25215 1285
rect 25285 1265 25300 1285
rect 25200 1250 25300 1265
rect 27200 1285 27300 1300
rect 27200 1265 27215 1285
rect 27285 1265 27300 1285
rect 27200 1250 27300 1265
rect 29200 1285 29300 1300
rect 29200 1265 29215 1285
rect 29285 1265 29300 1285
rect 29200 1250 29300 1265
rect 31200 1285 31300 1300
rect 31200 1265 31215 1285
rect 31285 1265 31300 1285
rect 31200 1250 31300 1265
rect 33200 1285 33300 1300
rect 33200 1265 33215 1285
rect 33285 1265 33300 1285
rect 33200 1250 33300 1265
rect 35200 1285 35300 1300
rect 35200 1265 35215 1285
rect 35285 1265 35300 1285
rect 35200 1250 35300 1265
rect 37200 1285 37300 1300
rect 37200 1265 37215 1285
rect 37285 1265 37300 1285
rect 37200 1250 37300 1265
rect 39200 1285 39300 1300
rect 39200 1265 39215 1285
rect 39285 1265 39300 1285
rect 39200 1250 39300 1265
rect 41200 1285 41300 1300
rect 41200 1265 41215 1285
rect 41285 1265 41300 1285
rect 41200 1250 41300 1265
rect 43200 1285 43300 1300
rect 43200 1265 43215 1285
rect 43285 1265 43300 1285
rect 43200 1250 43300 1265
rect 45200 1285 45300 1300
rect 45200 1265 45215 1285
rect 45285 1265 45300 1285
rect 45200 1250 45300 1265
rect 47200 1285 47300 1300
rect 47200 1265 47215 1285
rect 47285 1265 47300 1285
rect 47200 1250 47300 1265
rect 49200 1285 49300 1300
rect 49200 1265 49215 1285
rect 49285 1265 49300 1285
rect 49200 1250 49300 1265
rect 53550 1285 53650 1300
rect 53550 1265 53565 1285
rect 53635 1265 53650 1285
rect 53550 1250 53650 1265
rect 57550 1285 57650 1300
rect 57550 1265 57565 1285
rect 57635 1265 57650 1285
rect 57550 1250 57650 1265
<< psubdiffcont >>
rect 3215 1265 3285 1285
rect 5215 1265 5285 1285
rect 7215 1265 7285 1285
rect 9215 1265 9285 1285
rect 11215 1265 11285 1285
rect 13215 1265 13285 1285
rect 15215 1265 15285 1285
rect 17215 1265 17285 1285
rect 19215 1265 19285 1285
rect 21215 1265 21285 1285
rect 23215 1265 23285 1285
rect 25215 1265 25285 1285
rect 27215 1265 27285 1285
rect 29215 1265 29285 1285
rect 31215 1265 31285 1285
rect 33215 1265 33285 1285
rect 35215 1265 35285 1285
rect 37215 1265 37285 1285
rect 39215 1265 39285 1285
rect 41215 1265 41285 1285
rect 43215 1265 43285 1285
rect 45215 1265 45285 1285
rect 47215 1265 47285 1285
rect 49215 1265 49285 1285
rect 53565 1265 53635 1285
rect 57565 1265 57635 1285
<< locali >>
rect 3205 1285 3295 1295
rect 3205 1265 3215 1285
rect 3285 1265 3295 1285
rect 3205 1255 3295 1265
rect 5205 1285 5295 1295
rect 5205 1265 5215 1285
rect 5285 1265 5295 1285
rect 5205 1255 5295 1265
rect 7205 1285 7295 1295
rect 7205 1265 7215 1285
rect 7285 1265 7295 1285
rect 7205 1255 7295 1265
rect 9205 1285 9295 1295
rect 9205 1265 9215 1285
rect 9285 1265 9295 1285
rect 9205 1255 9295 1265
rect 11205 1285 11295 1295
rect 11205 1265 11215 1285
rect 11285 1265 11295 1285
rect 11205 1255 11295 1265
rect 13205 1285 13295 1295
rect 13205 1265 13215 1285
rect 13285 1265 13295 1285
rect 13205 1255 13295 1265
rect 15205 1285 15295 1295
rect 15205 1265 15215 1285
rect 15285 1265 15295 1285
rect 15205 1255 15295 1265
rect 17205 1285 17295 1295
rect 17205 1265 17215 1285
rect 17285 1265 17295 1285
rect 17205 1255 17295 1265
rect 19205 1285 19295 1295
rect 19205 1265 19215 1285
rect 19285 1265 19295 1285
rect 19205 1255 19295 1265
rect 21205 1285 21295 1295
rect 21205 1265 21215 1285
rect 21285 1265 21295 1285
rect 21205 1255 21295 1265
rect 23205 1285 23295 1295
rect 23205 1265 23215 1285
rect 23285 1265 23295 1285
rect 23205 1255 23295 1265
rect 25205 1285 25295 1295
rect 25205 1265 25215 1285
rect 25285 1265 25295 1285
rect 25205 1255 25295 1265
rect 27205 1285 27295 1295
rect 27205 1265 27215 1285
rect 27285 1265 27295 1285
rect 27205 1255 27295 1265
rect 29205 1285 29295 1295
rect 29205 1265 29215 1285
rect 29285 1265 29295 1285
rect 29205 1255 29295 1265
rect 31205 1285 31295 1295
rect 31205 1265 31215 1285
rect 31285 1265 31295 1285
rect 31205 1255 31295 1265
rect 33205 1285 33295 1295
rect 33205 1265 33215 1285
rect 33285 1265 33295 1285
rect 33205 1255 33295 1265
rect 35205 1285 35295 1295
rect 35205 1265 35215 1285
rect 35285 1265 35295 1285
rect 35205 1255 35295 1265
rect 37205 1285 37295 1295
rect 37205 1265 37215 1285
rect 37285 1265 37295 1285
rect 37205 1255 37295 1265
rect 39205 1285 39295 1295
rect 39205 1265 39215 1285
rect 39285 1265 39295 1285
rect 39205 1255 39295 1265
rect 41205 1285 41295 1295
rect 41205 1265 41215 1285
rect 41285 1265 41295 1285
rect 41205 1255 41295 1265
rect 43205 1285 43295 1295
rect 43205 1265 43215 1285
rect 43285 1265 43295 1285
rect 43205 1255 43295 1265
rect 45205 1285 45295 1295
rect 45205 1265 45215 1285
rect 45285 1265 45295 1285
rect 45205 1255 45295 1265
rect 47205 1285 47295 1295
rect 47205 1265 47215 1285
rect 47285 1265 47295 1285
rect 47205 1255 47295 1265
rect 49205 1285 49295 1295
rect 49205 1265 49215 1285
rect 49285 1265 49295 1285
rect 49205 1255 49295 1265
rect 53555 1285 53645 1295
rect 53555 1265 53565 1285
rect 53635 1265 53645 1285
rect 53555 1255 53645 1265
rect 57555 1285 57645 1295
rect 57555 1265 57565 1285
rect 57635 1265 57645 1285
rect 57555 1255 57645 1265
rect 7015 40 7035 360
rect 7875 40 7895 375
rect 7015 20 7315 40
rect 7450 20 7895 40
rect 14245 40 14265 385
rect 15105 40 15125 360
rect 21475 40 21495 365
rect 22335 40 22355 360
rect 14245 20 14560 40
rect 14695 20 15130 40
rect 21475 20 21855 40
rect 21915 20 22355 40
rect 28705 40 28725 380
rect 29565 40 29585 365
rect 28705 20 29045 40
rect 29180 20 29585 40
rect 35935 40 35955 370
rect 36795 40 36815 365
rect 35935 20 36315 40
rect 36410 20 36815 40
rect 43165 40 43185 360
rect 44025 40 44045 365
rect 43165 20 43575 40
rect 43680 20 44045 40
rect 50395 40 50415 360
rect 51255 40 51275 360
rect 50395 20 50770 40
rect 50905 20 51275 40
<< metal1 >>
rect 7230 215 58525 305
rect 7235 60 58525 145
use fvf  fvf_0
timestamp 1700263747
transform 1 0 39675 0 1 430
box -1790 1030 18445 8265
use inverter  inverter_0
timestamp 1693780072
transform 1 0 50980 0 1 145
box -240 -145 -30 185
use inverter  inverter_1
timestamp 1693780072
transform 1 0 7480 0 1 145
box -240 -145 -30 185
use inverter  inverter_2
timestamp 1693780072
transform 1 0 14730 0 1 145
box -240 -145 -30 185
use inverter  inverter_3
timestamp 1693780072
transform 1 0 21980 0 1 145
box -240 -145 -30 185
use inverter  inverter_4
timestamp 1693780072
transform 1 0 29230 0 1 145
box -240 -145 -30 185
use inverter  inverter_5
timestamp 1693780072
transform 1 0 36480 0 1 145
box -240 -145 -30 185
use inverter  inverter_6
timestamp 1693780072
transform 1 0 43730 0 1 145
box -240 -145 -30 185
use ladder  ladder_0
timestamp 1700206437
transform 1 0 10310 0 1 985
box -10460 -640 48210 205
<< end >>
