magic
tech sky130A
timestamp 1700322215
<< nmos >>
rect -8830 0 -8030 50
rect -7230 0 -6430 50
rect -5630 0 -4830 50
rect -4030 0 -3230 50
rect -2430 0 -1630 50
rect 0 0 800 50
rect 1600 0 2400 50
rect 3200 0 4000 50
rect 4800 0 5600 50
rect 7230 0 8030 50
rect 8830 0 9630 50
rect 10430 0 11230 50
rect 12030 0 12830 50
rect 14460 0 15260 50
rect 16060 0 16860 50
rect 17660 0 18460 50
rect 19260 0 20060 50
rect 21690 0 22490 50
rect 23290 0 24090 50
rect 24890 0 25690 50
rect 26490 0 27290 50
rect 28920 0 29720 50
rect 30520 0 31320 50
rect 32120 0 32920 50
rect 33720 0 34520 50
rect 36150 0 36950 50
rect 37750 0 38550 50
rect 39350 0 40150 50
rect 40950 0 41750 50
rect 43380 0 44180 50
rect 44980 0 45780 50
rect 46580 0 47380 50
rect -8830 -310 -8030 -260
rect -7230 -310 -6430 -260
rect -5630 -310 -4830 -260
rect -4030 -310 -3230 -260
rect -2430 -310 -1630 -260
rect 0 -310 800 -260
rect 1600 -310 2400 -260
rect 3200 -310 4000 -260
rect 4800 -310 5600 -260
rect 7230 -310 8030 -260
rect 8830 -310 9630 -260
rect 10430 -310 11230 -260
rect 12030 -310 12830 -260
rect 14460 -310 15260 -260
rect 16060 -310 16860 -260
rect 17660 -310 18460 -260
rect 19260 -310 20060 -260
rect 21690 -310 22490 -260
rect 23290 -310 24090 -260
rect 24890 -310 25690 -260
rect 26490 -310 27290 -260
rect 28920 -310 29720 -260
rect 30520 -310 31320 -260
rect 32120 -310 32920 -260
rect 33720 -310 34520 -260
rect 36150 -310 36950 -260
rect 37750 -310 38550 -260
rect 39350 -310 40150 -260
rect 40950 -310 41750 -260
rect 42550 -310 43350 -260
<< ndiff >>
rect -9630 35 -8830 50
rect -9630 15 -9615 35
rect -8845 15 -8830 35
rect -9630 0 -8830 15
rect -8030 35 -7230 50
rect -8030 15 -8015 35
rect -7245 15 -7230 35
rect -8030 0 -7230 15
rect -6430 35 -5630 50
rect -6430 15 -6415 35
rect -5645 15 -5630 35
rect -6430 0 -5630 15
rect -4830 35 -4030 50
rect -4830 15 -4815 35
rect -4045 15 -4030 35
rect -4830 0 -4030 15
rect -3230 35 -2430 50
rect -3230 15 -3215 35
rect -2445 15 -2430 35
rect -3230 0 -2430 15
rect -1630 35 -830 50
rect -1630 15 -1615 35
rect -845 15 -830 35
rect -1630 0 -830 15
rect -800 35 0 50
rect -800 15 -785 35
rect -15 15 0 35
rect -800 0 0 15
rect 800 35 1600 50
rect 800 15 815 35
rect 1585 15 1600 35
rect 800 0 1600 15
rect 2400 35 3200 50
rect 2400 15 2415 35
rect 3185 15 3200 35
rect 2400 0 3200 15
rect 4000 35 4800 50
rect 4000 15 4015 35
rect 4785 15 4800 35
rect 4000 0 4800 15
rect 5600 35 6400 50
rect 5600 15 5615 35
rect 6385 15 6400 35
rect 5600 0 6400 15
rect 6430 35 7230 50
rect 6430 15 6445 35
rect 7215 15 7230 35
rect 6430 0 7230 15
rect 8030 35 8830 50
rect 8030 15 8045 35
rect 8815 15 8830 35
rect 8030 0 8830 15
rect 9630 35 10430 50
rect 9630 15 9645 35
rect 10415 15 10430 35
rect 9630 0 10430 15
rect 11230 35 12030 50
rect 11230 15 11245 35
rect 12015 15 12030 35
rect 11230 0 12030 15
rect 12830 35 13630 50
rect 12830 15 12845 35
rect 13615 15 13630 35
rect 12830 0 13630 15
rect 13660 35 14460 50
rect 13660 15 13675 35
rect 14445 15 14460 35
rect 13660 0 14460 15
rect 15260 35 16060 50
rect 15260 15 15275 35
rect 16045 15 16060 35
rect 15260 0 16060 15
rect 16860 35 17660 50
rect 16860 15 16875 35
rect 17645 15 17660 35
rect 16860 0 17660 15
rect 18460 35 19260 50
rect 18460 15 18475 35
rect 19245 15 19260 35
rect 18460 0 19260 15
rect 20060 35 20860 50
rect 20060 15 20075 35
rect 20845 15 20860 35
rect 20060 0 20860 15
rect 20890 35 21690 50
rect 20890 15 20905 35
rect 21675 15 21690 35
rect 20890 0 21690 15
rect 22490 35 23290 50
rect 22490 15 22505 35
rect 23275 15 23290 35
rect 22490 0 23290 15
rect 24090 35 24890 50
rect 24090 15 24105 35
rect 24875 15 24890 35
rect 24090 0 24890 15
rect 25690 35 26490 50
rect 25690 15 25705 35
rect 26475 15 26490 35
rect 25690 0 26490 15
rect 27290 35 28090 50
rect 27290 15 27305 35
rect 28075 15 28090 35
rect 27290 0 28090 15
rect 28120 35 28920 50
rect 28120 15 28135 35
rect 28905 15 28920 35
rect 28120 0 28920 15
rect 29720 35 30520 50
rect 29720 15 29735 35
rect 30505 15 30520 35
rect 29720 0 30520 15
rect 31320 35 32120 50
rect 31320 15 31335 35
rect 32105 15 32120 35
rect 31320 0 32120 15
rect 32920 35 33720 50
rect 32920 15 32935 35
rect 33705 15 33720 35
rect 32920 0 33720 15
rect 34520 35 35320 50
rect 34520 15 34535 35
rect 35305 15 35320 35
rect 34520 0 35320 15
rect 35350 35 36150 50
rect 35350 15 35365 35
rect 36135 15 36150 35
rect 35350 0 36150 15
rect 36950 35 37750 50
rect 36950 15 36965 35
rect 37735 15 37750 35
rect 36950 0 37750 15
rect 38550 35 39350 50
rect 38550 15 38565 35
rect 39335 15 39350 35
rect 38550 0 39350 15
rect 40150 35 40950 50
rect 40150 15 40165 35
rect 40935 15 40950 35
rect 40150 0 40950 15
rect 41750 35 42550 50
rect 41750 15 41765 35
rect 42535 15 42550 35
rect 41750 0 42550 15
rect 42580 35 43380 50
rect 42580 15 42595 35
rect 43365 15 43380 35
rect 42580 0 43380 15
rect 44180 35 44980 50
rect 44180 15 44195 35
rect 44965 15 44980 35
rect 44180 0 44980 15
rect 45780 35 46580 50
rect 45780 15 45795 35
rect 46565 15 46580 35
rect 45780 0 46580 15
rect 47380 35 48180 50
rect 47380 15 47395 35
rect 48165 15 48180 35
rect 47380 0 48180 15
rect -9630 -275 -8830 -260
rect -9630 -295 -9615 -275
rect -8845 -295 -8830 -275
rect -9630 -310 -8830 -295
rect -8030 -275 -7230 -260
rect -8030 -295 -8015 -275
rect -7245 -295 -7230 -275
rect -8030 -310 -7230 -295
rect -6430 -275 -5630 -260
rect -6430 -295 -6415 -275
rect -5645 -295 -5630 -275
rect -6430 -310 -5630 -295
rect -4830 -275 -4030 -260
rect -4830 -295 -4815 -275
rect -4045 -295 -4030 -275
rect -4830 -310 -4030 -295
rect -3230 -275 -2430 -260
rect -3230 -295 -3215 -275
rect -2445 -295 -2430 -275
rect -3230 -310 -2430 -295
rect -1630 -275 -830 -260
rect -1630 -295 -1615 -275
rect -845 -295 -830 -275
rect -1630 -310 -830 -295
rect -800 -275 0 -260
rect -800 -295 -785 -275
rect -15 -295 0 -275
rect -800 -310 0 -295
rect 800 -275 1600 -260
rect 800 -295 815 -275
rect 1585 -295 1600 -275
rect 800 -310 1600 -295
rect 2400 -275 3200 -260
rect 2400 -295 2415 -275
rect 3185 -295 3200 -275
rect 2400 -310 3200 -295
rect 4000 -275 4800 -260
rect 4000 -295 4015 -275
rect 4785 -295 4800 -275
rect 4000 -310 4800 -295
rect 5600 -275 6400 -260
rect 5600 -295 5615 -275
rect 6385 -295 6400 -275
rect 5600 -310 6400 -295
rect 6430 -275 7230 -260
rect 6430 -295 6445 -275
rect 7215 -295 7230 -275
rect 6430 -310 7230 -295
rect 8030 -275 8830 -260
rect 8030 -295 8045 -275
rect 8815 -295 8830 -275
rect 8030 -310 8830 -295
rect 9630 -275 10430 -260
rect 9630 -295 9645 -275
rect 10415 -295 10430 -275
rect 9630 -310 10430 -295
rect 11230 -275 12030 -260
rect 11230 -295 11245 -275
rect 12015 -295 12030 -275
rect 11230 -310 12030 -295
rect 12830 -275 13630 -260
rect 12830 -295 12845 -275
rect 13615 -295 13630 -275
rect 12830 -310 13630 -295
rect 13660 -275 14460 -260
rect 13660 -295 13675 -275
rect 14445 -295 14460 -275
rect 13660 -310 14460 -295
rect 15260 -275 16060 -260
rect 15260 -295 15275 -275
rect 16045 -295 16060 -275
rect 15260 -310 16060 -295
rect 16860 -275 17660 -260
rect 16860 -295 16875 -275
rect 17645 -295 17660 -275
rect 16860 -310 17660 -295
rect 18460 -275 19260 -260
rect 18460 -295 18475 -275
rect 19245 -295 19260 -275
rect 18460 -310 19260 -295
rect 20060 -275 20860 -260
rect 20060 -295 20075 -275
rect 20845 -295 20860 -275
rect 20060 -310 20860 -295
rect 20890 -275 21690 -260
rect 20890 -295 20905 -275
rect 21675 -295 21690 -275
rect 20890 -310 21690 -295
rect 22490 -275 23290 -260
rect 22490 -295 22505 -275
rect 23275 -295 23290 -275
rect 22490 -310 23290 -295
rect 24090 -275 24890 -260
rect 24090 -295 24105 -275
rect 24875 -295 24890 -275
rect 24090 -310 24890 -295
rect 25690 -275 26490 -260
rect 25690 -295 25705 -275
rect 26475 -295 26490 -275
rect 25690 -310 26490 -295
rect 27290 -275 28090 -260
rect 27290 -295 27305 -275
rect 28075 -295 28090 -275
rect 27290 -310 28090 -295
rect 28120 -275 28920 -260
rect 28120 -295 28135 -275
rect 28905 -295 28920 -275
rect 28120 -310 28920 -295
rect 29720 -275 30520 -260
rect 29720 -295 29735 -275
rect 30505 -295 30520 -275
rect 29720 -310 30520 -295
rect 31320 -275 32120 -260
rect 31320 -295 31335 -275
rect 32105 -295 32120 -275
rect 31320 -310 32120 -295
rect 32920 -275 33720 -260
rect 32920 -295 32935 -275
rect 33705 -295 33720 -275
rect 32920 -310 33720 -295
rect 34520 -275 35320 -260
rect 34520 -295 34535 -275
rect 35305 -295 35320 -275
rect 34520 -310 35320 -295
rect 35350 -275 36150 -260
rect 35350 -295 35365 -275
rect 36135 -295 36150 -275
rect 35350 -310 36150 -295
rect 36950 -275 37750 -260
rect 36950 -295 36965 -275
rect 37735 -295 37750 -275
rect 36950 -310 37750 -295
rect 38550 -275 39350 -260
rect 38550 -295 38565 -275
rect 39335 -295 39350 -275
rect 38550 -310 39350 -295
rect 40150 -275 40950 -260
rect 40150 -295 40165 -275
rect 40935 -295 40950 -275
rect 40150 -310 40950 -295
rect 41750 -275 42550 -260
rect 41750 -295 41765 -275
rect 42535 -295 42550 -275
rect 41750 -310 42550 -295
rect 43350 -275 44150 -260
rect 43350 -295 43365 -275
rect 44135 -295 44150 -275
rect 43350 -310 44150 -295
<< ndiffc >>
rect -9615 15 -8845 35
rect -8015 15 -7245 35
rect -6415 15 -5645 35
rect -4815 15 -4045 35
rect -3215 15 -2445 35
rect -1615 15 -845 35
rect -785 15 -15 35
rect 815 15 1585 35
rect 2415 15 3185 35
rect 4015 15 4785 35
rect 5615 15 6385 35
rect 6445 15 7215 35
rect 8045 15 8815 35
rect 9645 15 10415 35
rect 11245 15 12015 35
rect 12845 15 13615 35
rect 13675 15 14445 35
rect 15275 15 16045 35
rect 16875 15 17645 35
rect 18475 15 19245 35
rect 20075 15 20845 35
rect 20905 15 21675 35
rect 22505 15 23275 35
rect 24105 15 24875 35
rect 25705 15 26475 35
rect 27305 15 28075 35
rect 28135 15 28905 35
rect 29735 15 30505 35
rect 31335 15 32105 35
rect 32935 15 33705 35
rect 34535 15 35305 35
rect 35365 15 36135 35
rect 36965 15 37735 35
rect 38565 15 39335 35
rect 40165 15 40935 35
rect 41765 15 42535 35
rect 42595 15 43365 35
rect 44195 15 44965 35
rect 45795 15 46565 35
rect 47395 15 48165 35
rect -9615 -295 -8845 -275
rect -8015 -295 -7245 -275
rect -6415 -295 -5645 -275
rect -4815 -295 -4045 -275
rect -3215 -295 -2445 -275
rect -1615 -295 -845 -275
rect -785 -295 -15 -275
rect 815 -295 1585 -275
rect 2415 -295 3185 -275
rect 4015 -295 4785 -275
rect 5615 -295 6385 -275
rect 6445 -295 7215 -275
rect 8045 -295 8815 -275
rect 9645 -295 10415 -275
rect 11245 -295 12015 -275
rect 12845 -295 13615 -275
rect 13675 -295 14445 -275
rect 15275 -295 16045 -275
rect 16875 -295 17645 -275
rect 18475 -295 19245 -275
rect 20075 -295 20845 -275
rect 20905 -295 21675 -275
rect 22505 -295 23275 -275
rect 24105 -295 24875 -275
rect 25705 -295 26475 -275
rect 27305 -295 28075 -275
rect 28135 -295 28905 -275
rect 29735 -295 30505 -275
rect 31335 -295 32105 -275
rect 32935 -295 33705 -275
rect 34535 -295 35305 -275
rect 35365 -295 36135 -275
rect 36965 -295 37735 -275
rect 38565 -295 39335 -275
rect 40165 -295 40935 -275
rect 41765 -295 42535 -275
rect 43365 -295 44135 -275
<< psubdiff >>
rect -7840 275 -7680 285
rect -7840 250 -7815 275
rect -7710 250 -7680 275
rect -7840 235 -7680 250
rect -5340 275 -5180 285
rect -5340 250 -5315 275
rect -5210 250 -5180 275
rect -5340 235 -5180 250
rect -2840 275 -2680 285
rect -2840 250 -2815 275
rect -2710 250 -2680 275
rect -2840 235 -2680 250
rect -340 275 -180 285
rect -340 250 -315 275
rect -210 250 -180 275
rect -340 235 -180 250
rect 2160 275 2320 285
rect 2160 250 2185 275
rect 2290 250 2320 275
rect 2160 235 2320 250
rect 4660 275 4820 285
rect 4660 250 4685 275
rect 4790 250 4820 275
rect 4660 235 4820 250
rect 7160 275 7320 285
rect 7160 250 7185 275
rect 7290 250 7320 275
rect 7160 235 7320 250
rect 9660 275 9820 285
rect 9660 250 9685 275
rect 9790 250 9820 275
rect 9660 235 9820 250
rect 12160 275 12320 285
rect 12160 250 12185 275
rect 12290 250 12320 275
rect 12160 235 12320 250
rect 14660 275 14820 285
rect 14660 250 14685 275
rect 14790 250 14820 275
rect 14660 235 14820 250
rect 17160 275 17320 285
rect 17160 250 17185 275
rect 17290 250 17320 275
rect 17160 235 17320 250
rect 19660 275 19820 285
rect 19660 250 19685 275
rect 19790 250 19820 275
rect 19660 235 19820 250
rect 22160 275 22320 285
rect 22160 250 22185 275
rect 22290 250 22320 275
rect 22160 235 22320 250
rect 24660 275 24820 285
rect 24660 250 24685 275
rect 24790 250 24820 275
rect 24660 235 24820 250
rect 27160 275 27320 285
rect 27160 250 27185 275
rect 27290 250 27320 275
rect 27160 235 27320 250
rect 29660 275 29820 285
rect 29660 250 29685 275
rect 29790 250 29820 275
rect 29660 235 29820 250
rect 32160 275 32320 285
rect 32160 250 32185 275
rect 32290 250 32320 275
rect 32160 235 32320 250
rect 34660 275 34820 285
rect 34660 250 34685 275
rect 34790 250 34820 275
rect 34660 235 34820 250
rect 37160 275 37320 285
rect 37160 250 37185 275
rect 37290 250 37320 275
rect 37160 235 37320 250
rect 39660 275 39820 285
rect 39660 250 39685 275
rect 39790 250 39820 275
rect 39660 235 39820 250
rect 42160 275 42320 285
rect 42160 250 42185 275
rect 42290 250 42320 275
rect 42160 235 42320 250
rect 44660 275 44820 285
rect 44660 250 44685 275
rect 44790 250 44820 275
rect 44660 235 44820 250
rect 47160 275 47320 285
rect 47160 250 47185 275
rect 47290 250 47320 275
rect 47160 235 47320 250
rect -10430 35 -9630 50
rect -10430 15 -10415 35
rect -9645 15 -9630 35
rect -10430 0 -9630 15
rect -10430 -275 -9630 -260
rect -10430 -295 -10415 -275
rect -9645 -295 -9630 -275
rect -10430 -310 -9630 -295
rect 44150 -275 44950 -260
rect 44150 -295 44160 -275
rect 44930 -295 44950 -275
rect 44150 -310 44950 -295
<< psubdiffcont >>
rect -7815 250 -7710 275
rect -5315 250 -5210 275
rect -2815 250 -2710 275
rect -315 250 -210 275
rect 2185 250 2290 275
rect 4685 250 4790 275
rect 7185 250 7290 275
rect 9685 250 9790 275
rect 12185 250 12290 275
rect 14685 250 14790 275
rect 17185 250 17290 275
rect 19685 250 19790 275
rect 22185 250 22290 275
rect 24685 250 24790 275
rect 27185 250 27290 275
rect 29685 250 29790 275
rect 32185 250 32290 275
rect 34685 250 34790 275
rect 37185 250 37290 275
rect 39685 250 39790 275
rect 42185 250 42290 275
rect 44685 250 44790 275
rect 47185 250 47290 275
rect -10415 15 -9645 35
rect -10415 -295 -9645 -275
rect 44160 -295 44930 -275
<< poly >>
rect -6090 155 -6045 165
rect -6090 135 -6080 155
rect -6055 140 -6045 155
rect -5785 155 -5740 165
rect -5785 140 -5775 155
rect -6055 135 -5775 140
rect -5750 135 -5740 155
rect -6090 125 -5740 135
rect -2960 155 -2915 165
rect -2960 135 -2950 155
rect -2925 140 -2915 155
rect -2725 155 -2680 165
rect -2725 140 -2715 155
rect -2925 135 -2715 140
rect -2690 135 -2680 155
rect -2960 125 -2680 135
rect 1140 155 1185 165
rect 1140 135 1150 155
rect 1175 140 1185 155
rect 1445 155 1490 165
rect 1445 140 1455 155
rect 1175 135 1455 140
rect 1480 135 1490 155
rect 1140 125 1490 135
rect 4270 155 4315 165
rect 4270 135 4280 155
rect 4305 140 4315 155
rect 4505 155 4550 165
rect 4505 140 4515 155
rect 4305 135 4515 140
rect 4540 135 4550 155
rect 4270 125 4550 135
rect 8370 155 8415 165
rect 8370 135 8380 155
rect 8405 140 8415 155
rect 8675 155 8720 165
rect 8675 140 8685 155
rect 8405 135 8685 140
rect 8710 135 8720 155
rect 8370 125 8720 135
rect 11500 155 11545 165
rect 11500 135 11510 155
rect 11535 140 11545 155
rect 11735 155 11780 165
rect 11735 140 11745 155
rect 11535 135 11745 140
rect 11770 135 11780 155
rect 11500 125 11780 135
rect 15600 155 15645 165
rect 15600 135 15610 155
rect 15635 140 15645 155
rect 15905 155 15950 165
rect 15905 140 15915 155
rect 15635 135 15915 140
rect 15940 135 15950 155
rect 15600 125 15950 135
rect 18730 155 18775 165
rect 18730 135 18740 155
rect 18765 140 18775 155
rect 18965 155 19010 165
rect 18965 140 18975 155
rect 18765 135 18975 140
rect 19000 135 19010 155
rect 18730 125 19010 135
rect 22830 155 22875 165
rect 22830 135 22840 155
rect 22865 140 22875 155
rect 23135 155 23180 165
rect 23135 140 23145 155
rect 22865 135 23145 140
rect 23170 135 23180 155
rect 22830 125 23180 135
rect 25960 155 26005 165
rect 25960 135 25970 155
rect 25995 140 26005 155
rect 26195 155 26240 165
rect 26195 140 26205 155
rect 25995 135 26205 140
rect 26230 135 26240 155
rect 25960 125 26240 135
rect 30060 155 30105 165
rect 30060 135 30070 155
rect 30095 140 30105 155
rect 30365 155 30410 165
rect 30365 140 30375 155
rect 30095 135 30375 140
rect 30400 135 30410 155
rect 30060 125 30410 135
rect 33190 155 33235 165
rect 33190 135 33200 155
rect 33225 140 33235 155
rect 33425 155 33470 165
rect 33425 140 33435 155
rect 33225 135 33435 140
rect 33460 135 33470 155
rect 33190 125 33470 135
rect 37290 155 37335 165
rect 37290 135 37300 155
rect 37325 140 37335 155
rect 37595 155 37640 165
rect 37595 140 37605 155
rect 37325 135 37605 140
rect 37630 135 37640 155
rect 37290 125 37640 135
rect 40420 155 40465 165
rect 40420 135 40430 155
rect 40455 140 40465 155
rect 40655 155 40700 165
rect 40655 140 40665 155
rect 40455 135 40665 140
rect 40690 135 40700 155
rect 40420 125 40700 135
rect -6500 95 -6455 100
rect -6500 75 -6490 95
rect -6465 75 -6455 95
rect -6500 65 -6455 75
rect -4900 95 -4855 100
rect -4900 75 -4890 95
rect -4865 75 -4855 95
rect -4900 65 -4855 75
rect -3300 95 -3255 100
rect -3300 75 -3290 95
rect -3265 75 -3255 95
rect -3300 65 -3255 75
rect -1700 95 -1655 100
rect -1700 75 -1690 95
rect -1665 75 -1655 95
rect -1700 65 -1655 75
rect 730 95 775 100
rect 730 75 740 95
rect 765 75 775 95
rect 730 65 775 75
rect 2330 95 2375 100
rect 2330 75 2340 95
rect 2365 75 2375 95
rect 2330 65 2375 75
rect 3930 95 3975 100
rect 3930 75 3940 95
rect 3965 75 3975 95
rect 3930 65 3975 75
rect 5530 95 5575 100
rect 5530 75 5540 95
rect 5565 75 5575 95
rect 5530 65 5575 75
rect 7960 95 8005 100
rect 7960 75 7970 95
rect 7995 75 8005 95
rect 7960 65 8005 75
rect 9560 95 9605 100
rect 9560 75 9570 95
rect 9595 75 9605 95
rect 9560 65 9605 75
rect 11160 95 11205 100
rect 11160 75 11170 95
rect 11195 75 11205 95
rect 11160 65 11205 75
rect 12760 95 12805 100
rect 12760 75 12770 95
rect 12795 75 12805 95
rect 12760 65 12805 75
rect 15190 95 15235 100
rect 15190 75 15200 95
rect 15225 75 15235 95
rect 15190 65 15235 75
rect 16790 95 16835 100
rect 16790 75 16800 95
rect 16825 75 16835 95
rect 16790 65 16835 75
rect 18390 95 18435 100
rect 18390 75 18400 95
rect 18425 75 18435 95
rect 18390 65 18435 75
rect 19990 95 20035 100
rect 19990 75 20000 95
rect 20025 75 20035 95
rect 19990 65 20035 75
rect 22420 95 22465 100
rect 22420 75 22430 95
rect 22455 75 22465 95
rect 22420 65 22465 75
rect 24020 95 24065 100
rect 24020 75 24030 95
rect 24055 75 24065 95
rect 24020 65 24065 75
rect 25620 95 25665 100
rect 25620 75 25630 95
rect 25655 75 25665 95
rect 25620 65 25665 75
rect 27220 95 27265 100
rect 27220 75 27230 95
rect 27255 75 27265 95
rect 27220 65 27265 75
rect 29650 95 29695 100
rect 29650 75 29660 95
rect 29685 75 29695 95
rect 29650 65 29695 75
rect 31250 95 31295 100
rect 31250 75 31260 95
rect 31285 75 31295 95
rect 31250 65 31295 75
rect 32850 95 32895 100
rect 32850 75 32860 95
rect 32885 75 32895 95
rect 32850 65 32895 75
rect 34450 95 34495 100
rect 34450 75 34460 95
rect 34485 75 34495 95
rect 34450 65 34495 75
rect 36880 95 36925 100
rect 36880 75 36890 95
rect 36915 75 36925 95
rect 36880 65 36925 75
rect 38480 95 38525 100
rect 38480 75 38490 95
rect 38515 75 38525 95
rect 38480 65 38525 75
rect 40080 95 40125 100
rect 40080 75 40090 95
rect 40115 75 40125 95
rect 40080 65 40125 75
rect 41680 95 41725 100
rect 41680 75 41690 95
rect 41715 75 41725 95
rect 41680 65 41725 75
rect 44110 95 44155 100
rect 44110 75 44120 95
rect 44145 75 44155 95
rect 44110 65 44155 75
rect 45710 95 45755 100
rect 45710 75 45720 95
rect 45745 75 45755 95
rect 45710 65 45755 75
rect 47310 90 47355 100
rect 47310 70 47320 90
rect 47345 70 47355 90
rect 47310 65 47355 70
rect -8830 50 -8030 65
rect -7230 50 -6430 65
rect -5630 50 -4830 65
rect -4030 50 -3230 65
rect -2430 50 -1630 65
rect 0 50 800 65
rect 1600 50 2400 65
rect 3200 50 4000 65
rect 4800 50 5600 65
rect 7230 50 8030 65
rect 8830 50 9630 65
rect 10430 50 11230 65
rect 12030 50 12830 65
rect 14460 50 15260 65
rect 16060 50 16860 65
rect 17660 50 18460 65
rect 19260 50 20060 65
rect 21690 50 22490 65
rect 23290 50 24090 65
rect 24890 50 25690 65
rect 26490 50 27290 65
rect 28920 50 29720 65
rect 30520 50 31320 65
rect 32120 50 32920 65
rect 33720 50 34520 65
rect 36150 50 36950 65
rect 37750 50 38550 65
rect 39350 50 40150 65
rect 40950 50 41750 65
rect 43380 50 44180 65
rect 44980 50 45780 65
rect 46580 50 47380 65
rect -8830 -15 -8030 0
rect -7230 -15 -6430 0
rect -5630 -15 -4830 0
rect -4030 -15 -3230 0
rect -2430 -15 -1630 0
rect 0 -15 800 0
rect 1600 -15 2400 0
rect 3200 -15 4000 0
rect 4800 -15 5600 0
rect 7230 -15 8030 0
rect 8830 -15 9630 0
rect 10430 -15 11230 0
rect 12030 -15 12830 0
rect 14460 -15 15260 0
rect 16060 -15 16860 0
rect 17660 -15 18460 0
rect 19260 -15 20060 0
rect 21690 -15 22490 0
rect 23290 -15 24090 0
rect 24890 -15 25690 0
rect 26490 -15 27290 0
rect 28920 -15 29720 0
rect 30520 -15 31320 0
rect 32120 -15 32920 0
rect 33720 -15 34520 0
rect 36150 -15 36950 0
rect 37750 -15 38550 0
rect 39350 -15 40150 0
rect 40950 -15 41750 0
rect 43380 -15 44180 0
rect 44980 -15 45780 0
rect 46580 -15 47380 0
rect -8805 -20 -8760 -15
rect -8805 -40 -8795 -20
rect -8770 -40 -8760 -20
rect -8805 -50 -8760 -40
rect -4530 -175 -4485 -165
rect -4530 -195 -4520 -175
rect -4495 -190 -4485 -175
rect -4365 -175 -4320 -165
rect -4365 -190 -4355 -175
rect -4495 -195 -4355 -190
rect -4330 -195 -4320 -175
rect -4530 -205 -4320 -195
rect 2700 -175 2745 -165
rect 2700 -195 2710 -175
rect 2735 -190 2745 -175
rect 2865 -175 2910 -165
rect 2865 -190 2875 -175
rect 2735 -195 2875 -190
rect 2900 -195 2910 -175
rect 2700 -205 2910 -195
rect 9930 -175 9975 -165
rect 9930 -195 9940 -175
rect 9965 -190 9975 -175
rect 10095 -175 10140 -165
rect 10095 -190 10105 -175
rect 9965 -195 10105 -190
rect 10130 -195 10140 -175
rect 9930 -205 10140 -195
rect 17160 -175 17205 -165
rect 17160 -195 17170 -175
rect 17195 -190 17205 -175
rect 17325 -175 17370 -165
rect 17325 -190 17335 -175
rect 17195 -195 17335 -190
rect 17360 -195 17370 -175
rect 17160 -205 17370 -195
rect 24390 -175 24435 -165
rect 24390 -195 24400 -175
rect 24425 -190 24435 -175
rect 24555 -175 24600 -165
rect 24555 -190 24565 -175
rect 24425 -195 24565 -190
rect 24590 -195 24600 -175
rect 24390 -205 24600 -195
rect 31620 -175 31665 -165
rect 31620 -195 31630 -175
rect 31655 -190 31665 -175
rect 31785 -175 31830 -165
rect 31785 -190 31795 -175
rect 31655 -195 31795 -190
rect 31820 -195 31830 -175
rect 31620 -205 31830 -195
rect 38850 -175 38895 -165
rect 38850 -195 38860 -175
rect 38885 -190 38895 -175
rect 39015 -175 39060 -165
rect 39015 -190 39025 -175
rect 38885 -195 39025 -190
rect 39050 -195 39060 -175
rect 38850 -205 39060 -195
rect 43280 -220 43325 -210
rect 43280 -240 43290 -220
rect 43315 -240 43325 -220
rect 43280 -245 43325 -240
rect -8830 -260 -8030 -245
rect -7230 -260 -6430 -245
rect -5630 -260 -4830 -245
rect -4030 -260 -3230 -245
rect -2430 -260 -1630 -245
rect 0 -260 800 -245
rect 1600 -260 2400 -245
rect 3200 -260 4000 -245
rect 4800 -260 5600 -245
rect 7230 -260 8030 -245
rect 8830 -260 9630 -245
rect 10430 -260 11230 -245
rect 12030 -260 12830 -245
rect 14460 -260 15260 -245
rect 16060 -260 16860 -245
rect 17660 -260 18460 -245
rect 19260 -260 20060 -245
rect 21690 -260 22490 -245
rect 23290 -260 24090 -245
rect 24890 -260 25690 -245
rect 26490 -260 27290 -245
rect 28920 -260 29720 -245
rect 30520 -260 31320 -245
rect 32120 -260 32920 -245
rect 33720 -260 34520 -245
rect 36150 -260 36950 -245
rect 37750 -260 38550 -245
rect 39350 -260 40150 -245
rect 40950 -260 41750 -245
rect 42550 -260 43350 -245
rect -8830 -325 -8030 -310
rect -7230 -325 -6430 -310
rect -5630 -325 -4830 -310
rect -4030 -325 -3230 -310
rect -2430 -325 -1630 -310
rect 0 -325 800 -310
rect 1600 -325 2400 -310
rect 3200 -325 4000 -310
rect 4800 -325 5600 -310
rect 7230 -325 8030 -310
rect 8830 -325 9630 -310
rect 10430 -325 11230 -310
rect 12030 -325 12830 -310
rect 14460 -325 15260 -310
rect 16060 -325 16860 -310
rect 17660 -325 18460 -310
rect 19260 -325 20060 -310
rect 21690 -325 22490 -310
rect 23290 -325 24090 -310
rect 24890 -325 25690 -310
rect 26490 -325 27290 -310
rect 28920 -325 29720 -310
rect 30520 -325 31320 -310
rect 32120 -325 32920 -310
rect 33720 -325 34520 -310
rect 36150 -325 36950 -310
rect 37750 -325 38550 -310
rect 39350 -325 40150 -310
rect 40950 -325 41750 -310
rect 42550 -325 43350 -310
rect -8805 -330 -8760 -325
rect -8805 -350 -8795 -330
rect -8770 -350 -8760 -330
rect -8805 -360 -8760 -350
rect -6445 -385 -6430 -325
rect -4845 -340 -4015 -325
rect -3300 -330 -3255 -325
rect -3300 -350 -3290 -330
rect -3265 -350 -3255 -330
rect -3300 -360 -3255 -350
rect -2430 -385 -2415 -325
rect -6445 -400 -2415 -385
rect 785 -385 800 -325
rect 2385 -340 3215 -325
rect 3930 -330 3975 -325
rect 3930 -350 3940 -330
rect 3965 -350 3975 -330
rect 3930 -360 3975 -350
rect 4800 -385 4815 -325
rect 785 -400 4815 -385
rect 8015 -385 8030 -325
rect 9615 -340 10445 -325
rect 11160 -330 11205 -325
rect 11160 -350 11170 -330
rect 11195 -350 11205 -330
rect 11160 -360 11205 -350
rect 12030 -385 12045 -325
rect 8015 -400 12045 -385
rect 15245 -385 15260 -325
rect 16845 -340 17675 -325
rect 18390 -330 18435 -325
rect 18390 -350 18400 -330
rect 18425 -350 18435 -330
rect 18390 -360 18435 -350
rect 19260 -385 19275 -325
rect 15245 -400 19275 -385
rect 22475 -385 22490 -325
rect 24075 -340 24905 -325
rect 25620 -330 25665 -325
rect 25620 -350 25630 -330
rect 25655 -350 25665 -330
rect 25620 -360 25665 -350
rect 26490 -385 26505 -325
rect 22475 -400 26505 -385
rect 29705 -385 29720 -325
rect 31305 -340 32135 -325
rect 32850 -330 32895 -325
rect 32850 -350 32860 -330
rect 32885 -350 32895 -330
rect 32850 -360 32895 -350
rect 33720 -385 33735 -325
rect 29705 -400 33735 -385
rect 36935 -385 36950 -325
rect 38535 -340 39365 -325
rect 40080 -330 40125 -325
rect 40080 -350 40090 -330
rect 40115 -350 40125 -330
rect 40080 -360 40125 -350
rect 40950 -385 40965 -325
rect 36935 -400 40965 -385
rect -4080 -440 -4035 -435
rect -4080 -460 -4070 -440
rect -4045 -460 -4035 -440
rect -4080 -470 -4035 -460
rect -3300 -440 -3255 -435
rect -3300 -460 -3290 -440
rect -3265 -460 -3255 -440
rect -3300 -470 -3255 -460
rect -4050 -530 -4035 -470
rect -4080 -540 -4035 -530
rect -4080 -560 -4070 -540
rect -4045 -560 -4035 -540
rect -4080 -565 -4035 -560
rect -3270 -570 -3255 -470
rect -2430 -570 -2415 -400
rect 3150 -440 3195 -435
rect 3150 -460 3160 -440
rect 3185 -460 3195 -440
rect 3150 -470 3195 -460
rect 3930 -440 3975 -435
rect 3930 -460 3940 -440
rect 3965 -460 3975 -440
rect 3930 -470 3975 -460
rect 3180 -530 3195 -470
rect 3150 -540 3195 -530
rect 3150 -560 3160 -540
rect 3185 -560 3195 -540
rect 3150 -565 3195 -560
rect 3960 -570 3975 -470
rect 4800 -570 4815 -400
rect 10380 -440 10425 -435
rect 10380 -460 10390 -440
rect 10415 -460 10425 -440
rect 10380 -470 10425 -460
rect 11160 -440 11205 -435
rect 11160 -460 11170 -440
rect 11195 -460 11205 -440
rect 11160 -470 11205 -460
rect 10410 -530 10425 -470
rect 10380 -540 10425 -530
rect 10380 -560 10390 -540
rect 10415 -560 10425 -540
rect 10380 -565 10425 -560
rect 11190 -570 11205 -470
rect 12030 -570 12045 -400
rect 17610 -440 17655 -435
rect 17610 -460 17620 -440
rect 17645 -460 17655 -440
rect 17610 -470 17655 -460
rect 18390 -440 18435 -435
rect 18390 -460 18400 -440
rect 18425 -460 18435 -440
rect 18390 -470 18435 -460
rect 17640 -530 17655 -470
rect 17610 -540 17655 -530
rect 17610 -560 17620 -540
rect 17645 -560 17655 -540
rect 17610 -565 17655 -560
rect 18420 -570 18435 -470
rect 19260 -570 19275 -400
rect 24840 -440 24885 -435
rect 24840 -460 24850 -440
rect 24875 -460 24885 -440
rect 24840 -470 24885 -460
rect 25620 -440 25665 -435
rect 25620 -460 25630 -440
rect 25655 -460 25665 -440
rect 25620 -470 25665 -460
rect 24870 -530 24885 -470
rect 24840 -540 24885 -530
rect 24840 -560 24850 -540
rect 24875 -560 24885 -540
rect 24840 -565 24885 -560
rect 25650 -570 25665 -470
rect 26490 -570 26505 -400
rect 32070 -440 32115 -435
rect 32070 -460 32080 -440
rect 32105 -460 32115 -440
rect 32070 -470 32115 -460
rect 32850 -440 32895 -435
rect 32850 -460 32860 -440
rect 32885 -460 32895 -440
rect 32850 -470 32895 -460
rect 32100 -530 32115 -470
rect 32070 -540 32115 -530
rect 32070 -560 32080 -540
rect 32105 -560 32115 -540
rect 32070 -565 32115 -560
rect 32880 -570 32895 -470
rect 33720 -570 33735 -400
rect 39300 -440 39345 -435
rect 39300 -460 39310 -440
rect 39335 -460 39345 -440
rect 39300 -470 39345 -460
rect 40080 -440 40125 -435
rect 40080 -460 40090 -440
rect 40115 -460 40125 -440
rect 40080 -470 40125 -460
rect 39330 -530 39345 -470
rect 39300 -540 39345 -530
rect 39300 -560 39310 -540
rect 39335 -560 39345 -540
rect 39300 -565 39345 -560
rect 40110 -570 40125 -470
rect 40950 -570 40965 -400
rect -3300 -580 -3255 -570
rect -3300 -600 -3290 -580
rect -3265 -600 -3255 -580
rect -3300 -605 -3255 -600
rect -2460 -580 -2415 -570
rect -2460 -600 -2450 -580
rect -2425 -600 -2415 -580
rect -2460 -605 -2415 -600
rect 3930 -580 3975 -570
rect 3930 -600 3940 -580
rect 3965 -600 3975 -580
rect 3930 -605 3975 -600
rect 4770 -580 4815 -570
rect 4770 -600 4780 -580
rect 4805 -600 4815 -580
rect 4770 -605 4815 -600
rect 11160 -580 11205 -570
rect 11160 -600 11170 -580
rect 11195 -600 11205 -580
rect 11160 -605 11205 -600
rect 12000 -580 12045 -570
rect 12000 -600 12010 -580
rect 12035 -600 12045 -580
rect 12000 -605 12045 -600
rect 18390 -580 18435 -570
rect 18390 -600 18400 -580
rect 18425 -600 18435 -580
rect 18390 -605 18435 -600
rect 19230 -580 19275 -570
rect 19230 -600 19240 -580
rect 19265 -600 19275 -580
rect 19230 -605 19275 -600
rect 25620 -580 25665 -570
rect 25620 -600 25630 -580
rect 25655 -600 25665 -580
rect 25620 -605 25665 -600
rect 26460 -580 26505 -570
rect 26460 -600 26470 -580
rect 26495 -600 26505 -580
rect 26460 -605 26505 -600
rect 32850 -580 32895 -570
rect 32850 -600 32860 -580
rect 32885 -600 32895 -580
rect 32850 -605 32895 -600
rect 33690 -580 33735 -570
rect 33690 -600 33700 -580
rect 33725 -600 33735 -580
rect 33690 -605 33735 -600
rect 40080 -580 40125 -570
rect 40080 -600 40090 -580
rect 40115 -600 40125 -580
rect 40080 -605 40125 -600
rect 40920 -580 40965 -570
rect 40920 -600 40930 -580
rect 40955 -600 40965 -580
rect 40920 -605 40965 -600
<< polycont >>
rect -6080 135 -6055 155
rect -5775 135 -5750 155
rect -2950 135 -2925 155
rect -2715 135 -2690 155
rect 1150 135 1175 155
rect 1455 135 1480 155
rect 4280 135 4305 155
rect 4515 135 4540 155
rect 8380 135 8405 155
rect 8685 135 8710 155
rect 11510 135 11535 155
rect 11745 135 11770 155
rect 15610 135 15635 155
rect 15915 135 15940 155
rect 18740 135 18765 155
rect 18975 135 19000 155
rect 22840 135 22865 155
rect 23145 135 23170 155
rect 25970 135 25995 155
rect 26205 135 26230 155
rect 30070 135 30095 155
rect 30375 135 30400 155
rect 33200 135 33225 155
rect 33435 135 33460 155
rect 37300 135 37325 155
rect 37605 135 37630 155
rect 40430 135 40455 155
rect 40665 135 40690 155
rect -6490 75 -6465 95
rect -4890 75 -4865 95
rect -3290 75 -3265 95
rect -1690 75 -1665 95
rect 740 75 765 95
rect 2340 75 2365 95
rect 3940 75 3965 95
rect 5540 75 5565 95
rect 7970 75 7995 95
rect 9570 75 9595 95
rect 11170 75 11195 95
rect 12770 75 12795 95
rect 15200 75 15225 95
rect 16800 75 16825 95
rect 18400 75 18425 95
rect 20000 75 20025 95
rect 22430 75 22455 95
rect 24030 75 24055 95
rect 25630 75 25655 95
rect 27230 75 27255 95
rect 29660 75 29685 95
rect 31260 75 31285 95
rect 32860 75 32885 95
rect 34460 75 34485 95
rect 36890 75 36915 95
rect 38490 75 38515 95
rect 40090 75 40115 95
rect 41690 75 41715 95
rect 44120 75 44145 95
rect 45720 75 45745 95
rect 47320 70 47345 90
rect -8795 -40 -8770 -20
rect -4520 -195 -4495 -175
rect -4355 -195 -4330 -175
rect 2710 -195 2735 -175
rect 2875 -195 2900 -175
rect 9940 -195 9965 -175
rect 10105 -195 10130 -175
rect 17170 -195 17195 -175
rect 17335 -195 17360 -175
rect 24400 -195 24425 -175
rect 24565 -195 24590 -175
rect 31630 -195 31655 -175
rect 31795 -195 31820 -175
rect 38860 -195 38885 -175
rect 39025 -195 39050 -175
rect 43290 -240 43315 -220
rect -8795 -350 -8770 -330
rect -3290 -350 -3265 -330
rect 3940 -350 3965 -330
rect 11170 -350 11195 -330
rect 18400 -350 18425 -330
rect 25630 -350 25655 -330
rect 32860 -350 32885 -330
rect 40090 -350 40115 -330
rect -4070 -460 -4045 -440
rect -3290 -460 -3265 -440
rect -4070 -560 -4045 -540
rect 3160 -460 3185 -440
rect 3940 -460 3965 -440
rect 3160 -560 3185 -540
rect 10390 -460 10415 -440
rect 11170 -460 11195 -440
rect 10390 -560 10415 -540
rect 17620 -460 17645 -440
rect 18400 -460 18425 -440
rect 17620 -560 17645 -540
rect 24850 -460 24875 -440
rect 25630 -460 25655 -440
rect 24850 -560 24875 -540
rect 32080 -460 32105 -440
rect 32860 -460 32885 -440
rect 32080 -560 32105 -540
rect 39310 -460 39335 -440
rect 40090 -460 40115 -440
rect 39310 -560 39335 -540
rect -3290 -600 -3265 -580
rect -2450 -600 -2425 -580
rect 3940 -600 3965 -580
rect 4780 -600 4805 -580
rect 11170 -600 11195 -580
rect 12010 -600 12035 -580
rect 18400 -600 18425 -580
rect 19240 -600 19265 -580
rect 25630 -600 25655 -580
rect 26470 -600 26495 -580
rect 32860 -600 32885 -580
rect 33700 -600 33725 -580
rect 40090 -600 40115 -580
rect 40930 -600 40955 -580
<< locali >>
rect -7830 275 -7690 280
rect -7830 250 -7815 275
rect -7710 250 -7690 275
rect -7830 240 -7690 250
rect -5330 275 -5190 280
rect -5330 250 -5315 275
rect -5210 250 -5190 275
rect -5330 240 -5190 250
rect -2830 275 -2690 280
rect -2830 250 -2815 275
rect -2710 250 -2690 275
rect -2830 240 -2690 250
rect -330 275 -190 280
rect -330 250 -315 275
rect -210 250 -190 275
rect -330 240 -190 250
rect 2170 275 2310 280
rect 2170 250 2185 275
rect 2290 250 2310 275
rect 2170 240 2310 250
rect 4670 275 4810 280
rect 4670 250 4685 275
rect 4790 250 4810 275
rect 4670 240 4810 250
rect 7170 275 7310 280
rect 7170 250 7185 275
rect 7290 250 7310 275
rect 7170 240 7310 250
rect 9670 275 9810 280
rect 9670 250 9685 275
rect 9790 250 9810 275
rect 9670 240 9810 250
rect 12170 275 12310 280
rect 12170 250 12185 275
rect 12290 250 12310 275
rect 12170 240 12310 250
rect 14670 275 14810 280
rect 14670 250 14685 275
rect 14790 250 14810 275
rect 14670 240 14810 250
rect 17170 275 17310 280
rect 17170 250 17185 275
rect 17290 250 17310 275
rect 17170 240 17310 250
rect 19670 275 19810 280
rect 19670 250 19685 275
rect 19790 250 19810 275
rect 19670 240 19810 250
rect 22170 275 22310 280
rect 22170 250 22185 275
rect 22290 250 22310 275
rect 22170 240 22310 250
rect 24670 275 24810 280
rect 24670 250 24685 275
rect 24790 250 24810 275
rect 24670 240 24810 250
rect 27170 275 27310 280
rect 27170 250 27185 275
rect 27290 250 27310 275
rect 27170 240 27310 250
rect 29670 275 29810 280
rect 29670 250 29685 275
rect 29790 250 29810 275
rect 29670 240 29810 250
rect 32170 275 32310 280
rect 32170 250 32185 275
rect 32290 250 32310 275
rect 32170 240 32310 250
rect 34670 275 34810 280
rect 34670 250 34685 275
rect 34790 250 34810 275
rect 34670 240 34810 250
rect 37170 275 37310 280
rect 37170 250 37185 275
rect 37290 250 37310 275
rect 37170 240 37310 250
rect 39670 275 39810 280
rect 39670 250 39685 275
rect 39790 250 39810 275
rect 39670 240 39810 250
rect 42170 275 42310 280
rect 42170 250 42185 275
rect 42290 250 42310 275
rect 42170 240 42310 250
rect 44670 275 44810 280
rect 44670 250 44685 275
rect 44790 250 44810 275
rect 44670 240 44810 250
rect 47170 275 47310 280
rect 47170 250 47185 275
rect 47290 250 47310 275
rect 47170 240 47310 250
rect -10460 185 -2820 205
rect -6090 155 -6045 165
rect -6090 145 -6080 155
rect -7255 135 -6080 145
rect -6055 135 -6045 155
rect -7255 125 -6045 135
rect -7255 45 -7235 125
rect -6500 95 -6455 100
rect -6500 75 -6490 95
rect -6465 75 -6455 95
rect -6500 65 -6455 75
rect -5945 45 -5925 185
rect -5785 155 -5740 165
rect -5785 135 -5775 155
rect -5750 145 -5740 155
rect -2960 155 -2915 165
rect -2960 145 -2950 155
rect -5750 135 -2950 145
rect -2925 135 -2915 155
rect -5785 125 -2915 135
rect -4900 95 -4855 100
rect -4900 75 -4890 95
rect -4865 75 -4855 95
rect -4900 65 -4855 75
rect -4435 65 -4415 100
rect -3300 95 -3255 100
rect -3300 75 -3290 95
rect -3265 75 -3255 95
rect -3300 65 -3255 75
rect -2840 45 -2820 185
rect -855 185 4410 205
rect -2725 155 -2680 165
rect -2725 135 -2715 155
rect -2690 145 -2680 155
rect -855 145 -835 185
rect 1140 155 1185 165
rect 1140 145 1150 155
rect -2690 135 -835 145
rect -2725 125 -835 135
rect -1700 95 -1655 100
rect -1700 75 -1690 95
rect -1665 75 -1655 95
rect -1700 65 -1655 75
rect -855 45 -835 125
rect -25 135 1150 145
rect 1175 135 1185 155
rect -25 125 1185 135
rect -25 45 -5 125
rect 730 95 775 100
rect 730 75 740 95
rect 765 75 775 95
rect 730 65 775 75
rect 1285 45 1305 185
rect 1445 155 1490 165
rect 1445 135 1455 155
rect 1480 145 1490 155
rect 4270 155 4315 165
rect 4270 145 4280 155
rect 1480 135 4280 145
rect 4305 135 4315 155
rect 1445 125 4315 135
rect 2330 95 2375 100
rect 2330 75 2340 95
rect 2365 75 2375 95
rect 2330 65 2375 75
rect 2795 65 2815 100
rect 3930 95 3975 100
rect 3930 75 3940 95
rect 3965 75 3975 95
rect 3930 65 3975 75
rect 4390 45 4410 185
rect 6375 185 11640 205
rect 4505 155 4550 165
rect 4505 135 4515 155
rect 4540 145 4550 155
rect 6375 145 6395 185
rect 8370 155 8415 165
rect 8370 145 8380 155
rect 4540 135 6395 145
rect 4505 125 6395 135
rect 5530 95 5575 100
rect 5530 75 5540 95
rect 5565 75 5575 95
rect 5530 65 5575 75
rect 6375 45 6395 125
rect 7205 135 8380 145
rect 8405 135 8415 155
rect 7205 125 8415 135
rect 7205 45 7225 125
rect 7960 95 8005 100
rect 7960 75 7970 95
rect 7995 75 8005 95
rect 7960 65 8005 75
rect 8515 45 8535 185
rect 8675 155 8720 165
rect 8675 135 8685 155
rect 8710 145 8720 155
rect 11500 155 11545 165
rect 11500 145 11510 155
rect 8710 135 11510 145
rect 11535 135 11545 155
rect 8675 125 11545 135
rect 9560 95 9605 100
rect 9560 75 9570 95
rect 9595 75 9605 95
rect 9560 65 9605 75
rect 10025 65 10045 100
rect 11160 95 11205 100
rect 11160 75 11170 95
rect 11195 75 11205 95
rect 11160 65 11205 75
rect 11620 45 11640 185
rect 13605 185 18870 205
rect 11735 155 11780 165
rect 11735 135 11745 155
rect 11770 145 11780 155
rect 13605 145 13625 185
rect 15600 155 15645 165
rect 15600 145 15610 155
rect 11770 135 13625 145
rect 11735 125 13625 135
rect 12760 95 12805 100
rect 12760 75 12770 95
rect 12795 75 12805 95
rect 12760 65 12805 75
rect 13605 45 13625 125
rect 14435 135 15610 145
rect 15635 135 15645 155
rect 14435 125 15645 135
rect 14435 45 14455 125
rect 15190 95 15235 100
rect 15190 75 15200 95
rect 15225 75 15235 95
rect 15190 65 15235 75
rect 15745 45 15765 185
rect 15905 155 15950 165
rect 15905 135 15915 155
rect 15940 145 15950 155
rect 18730 155 18775 165
rect 18730 145 18740 155
rect 15940 135 18740 145
rect 18765 135 18775 155
rect 15905 125 18775 135
rect 16790 95 16835 100
rect 16790 75 16800 95
rect 16825 75 16835 95
rect 16790 65 16835 75
rect 17255 65 17275 100
rect 18390 95 18435 100
rect 18390 75 18400 95
rect 18425 75 18435 95
rect 18390 65 18435 75
rect 18850 45 18870 185
rect 20835 185 26100 205
rect 18965 155 19010 165
rect 18965 135 18975 155
rect 19000 145 19010 155
rect 20835 145 20855 185
rect 22830 155 22875 165
rect 22830 145 22840 155
rect 19000 135 20855 145
rect 18965 125 20855 135
rect 19990 95 20035 100
rect 19990 75 20000 95
rect 20025 75 20035 95
rect 19990 65 20035 75
rect 20835 45 20855 125
rect 21665 135 22840 145
rect 22865 135 22875 155
rect 21665 125 22875 135
rect 21665 45 21685 125
rect 22420 95 22465 100
rect 22420 75 22430 95
rect 22455 75 22465 95
rect 22420 65 22465 75
rect 22975 45 22995 185
rect 23135 155 23180 165
rect 23135 135 23145 155
rect 23170 145 23180 155
rect 25960 155 26005 165
rect 25960 145 25970 155
rect 23170 135 25970 145
rect 25995 135 26005 155
rect 23135 125 26005 135
rect 24020 95 24065 100
rect 24020 75 24030 95
rect 24055 75 24065 95
rect 24020 65 24065 75
rect 24485 65 24505 100
rect 25620 95 25665 100
rect 25620 75 25630 95
rect 25655 75 25665 95
rect 25620 65 25665 75
rect 26080 45 26100 185
rect 28065 185 33330 205
rect 26195 155 26240 165
rect 26195 135 26205 155
rect 26230 145 26240 155
rect 28065 145 28085 185
rect 30060 155 30105 165
rect 30060 145 30070 155
rect 26230 135 28085 145
rect 26195 125 28085 135
rect 27220 95 27265 100
rect 27220 75 27230 95
rect 27255 75 27265 95
rect 27220 65 27265 75
rect 28065 45 28085 125
rect 28895 135 30070 145
rect 30095 135 30105 155
rect 28895 125 30105 135
rect 28895 45 28915 125
rect 29650 95 29695 100
rect 29650 75 29660 95
rect 29685 75 29695 95
rect 29650 65 29695 75
rect 30205 45 30225 185
rect 30365 155 30410 165
rect 30365 135 30375 155
rect 30400 145 30410 155
rect 33190 155 33235 165
rect 33190 145 33200 155
rect 30400 135 33200 145
rect 33225 135 33235 155
rect 30365 125 33235 135
rect 31250 95 31295 100
rect 31250 75 31260 95
rect 31285 75 31295 95
rect 31250 65 31295 75
rect 31715 65 31735 100
rect 32850 95 32895 100
rect 32850 75 32860 95
rect 32885 75 32895 95
rect 32850 65 32895 75
rect 33310 45 33330 185
rect 35295 185 40560 205
rect 33425 155 33470 165
rect 33425 135 33435 155
rect 33460 145 33470 155
rect 35295 145 35315 185
rect 37290 155 37335 165
rect 37290 145 37300 155
rect 33460 135 35315 145
rect 33425 125 35315 135
rect 34450 95 34495 100
rect 34450 75 34460 95
rect 34485 75 34495 95
rect 34450 65 34495 75
rect 35295 45 35315 125
rect 36125 135 37300 145
rect 37325 135 37335 155
rect 36125 125 37335 135
rect 36125 45 36145 125
rect 36880 95 36925 100
rect 36880 75 36890 95
rect 36915 75 36925 95
rect 36880 65 36925 75
rect 37435 45 37455 185
rect 37595 155 37640 165
rect 37595 135 37605 155
rect 37630 145 37640 155
rect 40420 155 40465 165
rect 40420 145 40430 155
rect 37630 135 40430 145
rect 40455 135 40465 155
rect 37595 125 40465 135
rect 38480 95 38525 100
rect 38480 75 38490 95
rect 38515 75 38525 95
rect 38480 65 38525 75
rect 38945 65 38965 100
rect 40080 95 40125 100
rect 40080 75 40090 95
rect 40115 75 40125 95
rect 40080 65 40125 75
rect 40540 45 40560 185
rect 42525 185 44205 205
rect 40655 155 40700 165
rect 40655 135 40665 155
rect 40690 145 40700 155
rect 42525 145 42545 185
rect 40690 135 42545 145
rect 40655 125 42545 135
rect 41680 95 41725 100
rect 41680 75 41690 95
rect 41715 75 41725 95
rect 41680 65 41725 75
rect 42525 45 42545 125
rect 44110 95 44155 100
rect 44110 75 44120 95
rect 44145 75 44155 95
rect 44110 65 44155 75
rect 44185 45 44205 185
rect 45710 95 45755 100
rect 45710 75 45720 95
rect 45745 75 45755 95
rect 45710 65 45755 75
rect 47310 90 47355 100
rect 47310 70 47320 90
rect 47345 85 47355 90
rect 47345 70 47405 85
rect 47310 65 47405 70
rect 47385 45 47405 65
rect -10425 35 -8835 45
rect -10425 15 -10415 35
rect -9645 15 -9615 35
rect -8845 15 -8835 35
rect -10425 5 -8835 15
rect -8025 35 -7235 45
rect -8025 15 -8015 35
rect -7245 15 -7235 35
rect -8025 5 -7235 15
rect -6425 35 -5635 45
rect -6425 15 -6415 35
rect -5645 15 -5635 35
rect -6425 5 -5635 15
rect -4825 35 -4035 45
rect -4825 15 -4815 35
rect -4045 15 -4035 35
rect -4825 5 -4035 15
rect -3225 35 -2435 45
rect -3225 15 -3215 35
rect -2445 15 -2435 35
rect -3225 5 -2435 15
rect -1625 35 -835 45
rect -1625 15 -1615 35
rect -845 15 -835 35
rect -1625 5 -835 15
rect -795 35 -5 45
rect -795 15 -785 35
rect -15 15 -5 35
rect -795 5 -5 15
rect 805 35 1595 45
rect 805 15 815 35
rect 1585 15 1595 35
rect 805 5 1595 15
rect 2405 35 3195 45
rect 2405 15 2415 35
rect 3185 15 3195 35
rect 2405 5 3195 15
rect 4005 35 4795 45
rect 4005 15 4015 35
rect 4785 15 4795 35
rect 4005 5 4795 15
rect 5605 35 6395 45
rect 5605 15 5615 35
rect 6385 15 6395 35
rect 5605 5 6395 15
rect 6435 35 7225 45
rect 6435 15 6445 35
rect 7215 15 7225 35
rect 6435 5 7225 15
rect 8035 35 8825 45
rect 8035 15 8045 35
rect 8815 15 8825 35
rect 8035 5 8825 15
rect 9635 35 10425 45
rect 9635 15 9645 35
rect 10415 15 10425 35
rect 9635 5 10425 15
rect 11235 35 12025 45
rect 11235 15 11245 35
rect 12015 15 12025 35
rect 11235 5 12025 15
rect 12835 35 13625 45
rect 12835 15 12845 35
rect 13615 15 13625 35
rect 12835 5 13625 15
rect 13665 35 14455 45
rect 13665 15 13675 35
rect 14445 15 14455 35
rect 13665 5 14455 15
rect 15265 35 16055 45
rect 15265 15 15275 35
rect 16045 15 16055 35
rect 15265 5 16055 15
rect 16865 35 17655 45
rect 16865 15 16875 35
rect 17645 15 17655 35
rect 16865 5 17655 15
rect 18465 35 19255 45
rect 18465 15 18475 35
rect 19245 15 19255 35
rect 18465 5 19255 15
rect 20065 35 20855 45
rect 20065 15 20075 35
rect 20845 15 20855 35
rect 20065 5 20855 15
rect 20895 35 21685 45
rect 20895 15 20905 35
rect 21675 15 21685 35
rect 20895 5 21685 15
rect 22495 35 23285 45
rect 22495 15 22505 35
rect 23275 15 23285 35
rect 22495 5 23285 15
rect 24095 35 24885 45
rect 24095 15 24105 35
rect 24875 15 24885 35
rect 24095 5 24885 15
rect 25695 35 26485 45
rect 25695 15 25705 35
rect 26475 15 26485 35
rect 25695 5 26485 15
rect 27295 35 28085 45
rect 27295 15 27305 35
rect 28075 15 28085 35
rect 27295 5 28085 15
rect 28125 35 28915 45
rect 28125 15 28135 35
rect 28905 15 28915 35
rect 28125 5 28915 15
rect 29725 35 30515 45
rect 29725 15 29735 35
rect 30505 15 30515 35
rect 29725 5 30515 15
rect 31325 35 32115 45
rect 31325 15 31335 35
rect 32105 15 32115 35
rect 31325 5 32115 15
rect 32925 35 33715 45
rect 32925 15 32935 35
rect 33705 15 33715 35
rect 32925 5 33715 15
rect 34525 35 35315 45
rect 34525 15 34535 35
rect 35305 15 35315 35
rect 34525 5 35315 15
rect 35355 35 36145 45
rect 35355 15 35365 35
rect 36135 15 36145 35
rect 35355 5 36145 15
rect 36955 35 37745 45
rect 36955 15 36965 35
rect 37735 15 37745 35
rect 36955 5 37745 15
rect 38555 35 39345 45
rect 38555 15 38565 35
rect 39335 15 39345 35
rect 38555 5 39345 15
rect 40155 35 40945 45
rect 40155 15 40165 35
rect 40935 15 40945 35
rect 40155 5 40945 15
rect 41755 35 42545 45
rect 41755 15 41765 35
rect 42535 15 42545 35
rect 41755 5 42545 15
rect 42585 35 43375 45
rect 42585 15 42595 35
rect 43365 15 43375 35
rect 42585 5 43375 15
rect 44185 35 44975 45
rect 44185 15 44195 35
rect 44965 15 44975 35
rect 44185 5 44975 15
rect 45785 35 46575 45
rect 45785 15 45795 35
rect 46565 15 46575 35
rect 45785 5 46575 15
rect 47385 35 48175 45
rect 47385 15 47395 35
rect 48165 15 48175 35
rect 47385 5 48175 15
rect -8855 -15 -8835 5
rect -8855 -20 -8760 -15
rect -8855 -35 -8795 -20
rect -8805 -40 -8795 -35
rect -8770 -40 -8760 -20
rect -8805 -50 -8760 -40
rect -4530 -175 -4485 -165
rect -4530 -185 -4520 -175
rect -7255 -195 -4520 -185
rect -4495 -195 -4485 -175
rect -7255 -205 -4485 -195
rect -7255 -265 -7235 -205
rect -4435 -225 -4415 5
rect -4365 -175 -4320 -165
rect -4365 -195 -4355 -175
rect -4330 -185 -4320 -175
rect 2700 -175 2745 -165
rect 2700 -185 2710 -175
rect -4330 -195 -1605 -185
rect -4365 -205 -1605 -195
rect -5655 -245 -3205 -225
rect -5655 -265 -5635 -245
rect -3225 -265 -3205 -245
rect -1625 -265 -1605 -205
rect -25 -195 2710 -185
rect 2735 -195 2745 -175
rect -25 -205 2745 -195
rect -25 -265 -5 -205
rect 2795 -225 2815 5
rect 2865 -175 2910 -165
rect 2865 -195 2875 -175
rect 2900 -185 2910 -175
rect 9930 -175 9975 -165
rect 9930 -185 9940 -175
rect 2900 -195 5625 -185
rect 2865 -205 5625 -195
rect 1575 -245 4025 -225
rect 1575 -265 1595 -245
rect 4005 -265 4025 -245
rect 5605 -265 5625 -205
rect 7205 -195 9940 -185
rect 9965 -195 9975 -175
rect 7205 -205 9975 -195
rect 7205 -265 7225 -205
rect 10025 -225 10045 5
rect 10095 -175 10140 -165
rect 10095 -195 10105 -175
rect 10130 -185 10140 -175
rect 17160 -175 17205 -165
rect 17160 -185 17170 -175
rect 10130 -195 12855 -185
rect 10095 -205 12855 -195
rect 8805 -245 11255 -225
rect 8805 -265 8825 -245
rect 11235 -265 11255 -245
rect 12835 -265 12855 -205
rect 14435 -195 17170 -185
rect 17195 -195 17205 -175
rect 14435 -205 17205 -195
rect 14435 -265 14455 -205
rect 17255 -225 17275 5
rect 17325 -175 17370 -165
rect 17325 -195 17335 -175
rect 17360 -185 17370 -175
rect 24390 -175 24435 -165
rect 24390 -185 24400 -175
rect 17360 -195 20085 -185
rect 17325 -205 20085 -195
rect 16035 -245 18485 -225
rect 16035 -265 16055 -245
rect 18465 -265 18485 -245
rect 20065 -265 20085 -205
rect 21665 -195 24400 -185
rect 24425 -195 24435 -175
rect 21665 -205 24435 -195
rect 21665 -265 21685 -205
rect 24485 -225 24505 5
rect 24555 -175 24600 -165
rect 24555 -195 24565 -175
rect 24590 -185 24600 -175
rect 31620 -175 31665 -165
rect 31620 -185 31630 -175
rect 24590 -195 27315 -185
rect 24555 -205 27315 -195
rect 23265 -245 25715 -225
rect 23265 -265 23285 -245
rect 25695 -265 25715 -245
rect 27295 -265 27315 -205
rect 28895 -195 31630 -185
rect 31655 -195 31665 -175
rect 28895 -205 31665 -195
rect 28895 -265 28915 -205
rect 31715 -225 31735 5
rect 31785 -175 31830 -165
rect 31785 -195 31795 -175
rect 31820 -185 31830 -175
rect 38850 -175 38895 -165
rect 38850 -185 38860 -175
rect 31820 -195 34545 -185
rect 31785 -205 34545 -195
rect 30495 -245 32945 -225
rect 30495 -265 30515 -245
rect 32925 -265 32945 -245
rect 34525 -265 34545 -205
rect 36125 -195 38860 -185
rect 38885 -195 38895 -175
rect 36125 -205 38895 -195
rect 36125 -265 36145 -205
rect 38945 -225 38965 5
rect 43355 -15 43375 5
rect 45785 -15 45805 5
rect 43355 -35 45805 -15
rect 39015 -175 39060 -165
rect 39015 -195 39025 -175
rect 39050 -185 39060 -175
rect 39050 -195 41775 -185
rect 39015 -205 41775 -195
rect 37725 -245 40175 -225
rect 37725 -265 37745 -245
rect 40155 -265 40175 -245
rect 41755 -265 41775 -205
rect 43280 -220 43325 -210
rect 43280 -240 43290 -220
rect 43315 -240 43375 -220
rect 43280 -245 43325 -240
rect 43355 -265 43375 -240
rect -10425 -275 -8835 -265
rect -10425 -295 -10415 -275
rect -9645 -295 -9615 -275
rect -8845 -295 -8835 -275
rect -10425 -305 -8835 -295
rect -8025 -275 -7235 -265
rect -8025 -295 -8015 -275
rect -7245 -295 -7235 -275
rect -8025 -305 -7235 -295
rect -6425 -275 -5635 -265
rect -6425 -295 -6415 -275
rect -5645 -295 -5635 -275
rect -6425 -305 -5635 -295
rect -4825 -275 -4035 -265
rect -4825 -295 -4815 -275
rect -4045 -295 -4035 -275
rect -4825 -305 -4035 -295
rect -3225 -275 -2435 -265
rect -3225 -295 -3215 -275
rect -2445 -295 -2435 -275
rect -3225 -305 -2435 -295
rect -1625 -275 -835 -265
rect -1625 -295 -1615 -275
rect -845 -295 -835 -275
rect -1625 -305 -835 -295
rect -795 -275 -5 -265
rect -795 -295 -785 -275
rect -15 -295 -5 -275
rect -795 -305 -5 -295
rect 805 -275 1595 -265
rect 805 -295 815 -275
rect 1585 -295 1595 -275
rect 805 -305 1595 -295
rect 2405 -275 3195 -265
rect 2405 -295 2415 -275
rect 3185 -295 3195 -275
rect 2405 -305 3195 -295
rect 4005 -275 4795 -265
rect 4005 -295 4015 -275
rect 4785 -295 4795 -275
rect 4005 -305 4795 -295
rect 5605 -275 6395 -265
rect 5605 -295 5615 -275
rect 6385 -295 6395 -275
rect 5605 -305 6395 -295
rect 6435 -275 7225 -265
rect 6435 -295 6445 -275
rect 7215 -295 7225 -275
rect 6435 -305 7225 -295
rect 8035 -275 8825 -265
rect 8035 -295 8045 -275
rect 8815 -295 8825 -275
rect 8035 -305 8825 -295
rect 9635 -275 10425 -265
rect 9635 -295 9645 -275
rect 10415 -295 10425 -275
rect 9635 -305 10425 -295
rect 11235 -275 12025 -265
rect 11235 -295 11245 -275
rect 12015 -295 12025 -275
rect 11235 -305 12025 -295
rect 12835 -275 13625 -265
rect 12835 -295 12845 -275
rect 13615 -295 13625 -275
rect 12835 -305 13625 -295
rect 13665 -275 14455 -265
rect 13665 -295 13675 -275
rect 14445 -295 14455 -275
rect 13665 -305 14455 -295
rect 15265 -275 16055 -265
rect 15265 -295 15275 -275
rect 16045 -295 16055 -275
rect 15265 -305 16055 -295
rect 16865 -275 17655 -265
rect 16865 -295 16875 -275
rect 17645 -295 17655 -275
rect 16865 -305 17655 -295
rect 18465 -275 19255 -265
rect 18465 -295 18475 -275
rect 19245 -295 19255 -275
rect 18465 -305 19255 -295
rect 20065 -275 20855 -265
rect 20065 -295 20075 -275
rect 20845 -295 20855 -275
rect 20065 -305 20855 -295
rect 20895 -275 21685 -265
rect 20895 -295 20905 -275
rect 21675 -295 21685 -275
rect 20895 -305 21685 -295
rect 22495 -275 23285 -265
rect 22495 -295 22505 -275
rect 23275 -295 23285 -275
rect 22495 -305 23285 -295
rect 24095 -275 24885 -265
rect 24095 -295 24105 -275
rect 24875 -295 24885 -275
rect 24095 -305 24885 -295
rect 25695 -275 26485 -265
rect 25695 -295 25705 -275
rect 26475 -295 26485 -275
rect 25695 -305 26485 -295
rect 27295 -275 28085 -265
rect 27295 -295 27305 -275
rect 28075 -295 28085 -275
rect 27295 -305 28085 -295
rect 28125 -275 28915 -265
rect 28125 -295 28135 -275
rect 28905 -295 28915 -275
rect 28125 -305 28915 -295
rect 29725 -275 30515 -265
rect 29725 -295 29735 -275
rect 30505 -295 30515 -275
rect 29725 -305 30515 -295
rect 31325 -275 32115 -265
rect 31325 -295 31335 -275
rect 32105 -295 32115 -275
rect 31325 -305 32115 -295
rect 32925 -275 33715 -265
rect 32925 -295 32935 -275
rect 33705 -295 33715 -275
rect 32925 -305 33715 -295
rect 34525 -275 35315 -265
rect 34525 -295 34535 -275
rect 35305 -295 35315 -275
rect 34525 -305 35315 -295
rect 35355 -275 36145 -265
rect 35355 -295 35365 -275
rect 36135 -295 36145 -275
rect 35355 -305 36145 -295
rect 36955 -275 37745 -265
rect 36955 -295 36965 -275
rect 37735 -295 37745 -275
rect 36955 -305 37745 -295
rect 38555 -275 39345 -265
rect 38555 -295 38565 -275
rect 39335 -295 39345 -275
rect 38555 -305 39345 -295
rect 40155 -275 40945 -265
rect 40155 -295 40165 -275
rect 40935 -295 40945 -275
rect 40155 -305 40945 -295
rect 41755 -275 42545 -265
rect 41755 -295 41765 -275
rect 42535 -295 42545 -275
rect 41755 -305 42545 -295
rect 43355 -275 44945 -265
rect 43355 -295 43365 -275
rect 44135 -295 44160 -275
rect 44930 -295 44945 -275
rect 43355 -305 44945 -295
rect -8855 -325 -8835 -305
rect -8855 -330 -8760 -325
rect -8855 -345 -8795 -330
rect -8805 -350 -8795 -345
rect -8770 -350 -8760 -330
rect -8805 -360 -8760 -350
rect -4055 -435 -4035 -305
rect -3300 -330 -3255 -325
rect -3300 -350 -3290 -330
rect -3265 -350 -3255 -330
rect -3300 -360 -3255 -350
rect -3275 -435 -3255 -360
rect -4080 -440 -4035 -435
rect -4080 -460 -4070 -440
rect -4045 -460 -4035 -440
rect -4080 -470 -4035 -460
rect -3300 -440 -3255 -435
rect -3300 -460 -3290 -440
rect -3265 -460 -3255 -440
rect -3300 -470 -3255 -460
rect -855 -490 -835 -305
rect 3175 -435 3195 -305
rect 3930 -330 3975 -325
rect 3930 -350 3940 -330
rect 3965 -350 3975 -330
rect 3930 -360 3975 -350
rect 3955 -435 3975 -360
rect 3150 -440 3195 -435
rect 3150 -460 3160 -440
rect 3185 -460 3195 -440
rect 3150 -470 3195 -460
rect 3930 -440 3975 -435
rect 3930 -460 3940 -440
rect 3965 -460 3975 -440
rect 3930 -470 3975 -460
rect 6375 -490 6395 -305
rect 10405 -435 10425 -305
rect 11160 -330 11205 -325
rect 11160 -350 11170 -330
rect 11195 -350 11205 -330
rect 11160 -360 11205 -350
rect 11185 -435 11205 -360
rect 10380 -440 10425 -435
rect 10380 -460 10390 -440
rect 10415 -460 10425 -440
rect 10380 -470 10425 -460
rect 11160 -440 11205 -435
rect 11160 -460 11170 -440
rect 11195 -460 11205 -440
rect 11160 -470 11205 -460
rect 13605 -490 13625 -305
rect 17635 -435 17655 -305
rect 18390 -330 18435 -325
rect 18390 -350 18400 -330
rect 18425 -350 18435 -330
rect 18390 -360 18435 -350
rect 18415 -435 18435 -360
rect 17610 -440 17655 -435
rect 17610 -460 17620 -440
rect 17645 -460 17655 -440
rect 17610 -470 17655 -460
rect 18390 -440 18435 -435
rect 18390 -460 18400 -440
rect 18425 -460 18435 -440
rect 18390 -470 18435 -460
rect 20835 -490 20855 -305
rect 24865 -435 24885 -305
rect 25620 -330 25665 -325
rect 25620 -350 25630 -330
rect 25655 -350 25665 -330
rect 25620 -360 25665 -350
rect 25645 -435 25665 -360
rect 24840 -440 24885 -435
rect 24840 -460 24850 -440
rect 24875 -460 24885 -440
rect 24840 -470 24885 -460
rect 25620 -440 25665 -435
rect 25620 -460 25630 -440
rect 25655 -460 25665 -440
rect 25620 -470 25665 -460
rect 28065 -490 28085 -305
rect 32095 -435 32115 -305
rect 32850 -330 32895 -325
rect 32850 -350 32860 -330
rect 32885 -350 32895 -330
rect 32850 -360 32895 -350
rect 32875 -435 32895 -360
rect 32070 -440 32115 -435
rect 32070 -460 32080 -440
rect 32105 -460 32115 -440
rect 32070 -470 32115 -460
rect 32850 -440 32895 -435
rect 32850 -460 32860 -440
rect 32885 -460 32895 -440
rect 32850 -470 32895 -460
rect 35295 -490 35315 -305
rect 39325 -435 39345 -305
rect 40080 -330 40125 -325
rect 40080 -350 40090 -330
rect 40115 -350 40125 -330
rect 40080 -360 40125 -350
rect 40105 -435 40125 -360
rect 39300 -440 39345 -435
rect 39300 -460 39310 -440
rect 39335 -460 39345 -440
rect 39300 -470 39345 -460
rect 40080 -440 40125 -435
rect 40080 -460 40090 -440
rect 40115 -460 40125 -440
rect 40080 -470 40125 -460
rect 42525 -490 42545 -305
rect 45785 -490 45805 -35
rect -4080 -510 48210 -490
rect -4080 -540 48210 -530
rect -4080 -560 -4070 -540
rect -4045 -550 3160 -540
rect -4045 -560 -4035 -550
rect -4080 -565 -4035 -560
rect 3150 -560 3160 -550
rect 3185 -550 10390 -540
rect 3185 -560 3195 -550
rect 3150 -565 3195 -560
rect 10380 -560 10390 -550
rect 10415 -550 17620 -540
rect 10415 -560 10425 -550
rect 10380 -565 10425 -560
rect 17610 -560 17620 -550
rect 17645 -550 24850 -540
rect 17645 -560 17655 -550
rect 17610 -565 17655 -560
rect 24840 -560 24850 -550
rect 24875 -550 32080 -540
rect 24875 -560 24885 -550
rect 24840 -565 24885 -560
rect 32070 -560 32080 -550
rect 32105 -550 39310 -540
rect 32105 -560 32115 -550
rect 32070 -565 32115 -560
rect 39300 -560 39310 -550
rect 39335 -550 48210 -540
rect 39335 -560 39345 -550
rect 39300 -565 39345 -560
rect -3300 -580 -3255 -570
rect -3300 -600 -3290 -580
rect -3265 -600 -3255 -580
rect -3300 -605 -3255 -600
rect -2460 -580 -2415 -570
rect -2460 -600 -2450 -580
rect -2425 -600 -2415 -580
rect -2460 -605 -2415 -600
rect 3930 -580 3975 -570
rect 3930 -600 3940 -580
rect 3965 -600 3975 -580
rect 3930 -605 3975 -600
rect 4770 -580 4815 -570
rect 4770 -600 4780 -580
rect 4805 -600 4815 -580
rect 4770 -605 4815 -600
rect 11160 -580 11205 -570
rect 11160 -600 11170 -580
rect 11195 -600 11205 -580
rect 11160 -605 11205 -600
rect 12000 -580 12045 -570
rect 12000 -600 12010 -580
rect 12035 -600 12045 -580
rect 12000 -605 12045 -600
rect 18390 -580 18435 -570
rect 18390 -600 18400 -580
rect 18425 -600 18435 -580
rect 18390 -605 18435 -600
rect 19230 -580 19275 -570
rect 19230 -600 19240 -580
rect 19265 -600 19275 -580
rect 19230 -605 19275 -600
rect 25620 -580 25665 -570
rect 25620 -600 25630 -580
rect 25655 -600 25665 -580
rect 25620 -605 25665 -600
rect 26460 -580 26505 -570
rect 26460 -600 26470 -580
rect 26495 -600 26505 -580
rect 26460 -605 26505 -600
rect 32850 -580 32895 -570
rect 32850 -600 32860 -580
rect 32885 -600 32895 -580
rect 32850 -605 32895 -600
rect 33690 -580 33735 -570
rect 33690 -600 33700 -580
rect 33725 -600 33735 -580
rect 33690 -605 33735 -600
rect 40080 -580 40125 -570
rect 40080 -600 40090 -580
rect 40115 -600 40125 -580
rect 40080 -605 40125 -600
rect 40920 -580 40965 -570
rect 40920 -600 40930 -580
rect 40955 -600 40965 -580
rect 40920 -605 40965 -600
rect -3295 -640 -3275 -605
rect -2435 -640 -2415 -605
rect 3935 -640 3955 -605
rect 4795 -640 4815 -605
rect 11165 -640 11185 -605
rect 12025 -640 12045 -605
rect 18395 -640 18415 -605
rect 19255 -640 19275 -605
rect 25625 -640 25645 -605
rect 26485 -640 26505 -605
rect 32855 -640 32875 -605
rect 33715 -640 33735 -605
rect 40085 -640 40105 -605
rect 40945 -640 40965 -605
<< viali >>
rect -7815 250 -7710 275
rect -5315 250 -5210 275
rect -2815 250 -2710 275
rect -315 250 -210 275
rect 2185 250 2290 275
rect 4685 250 4790 275
rect 7185 250 7290 275
rect 9685 250 9790 275
rect 12185 250 12290 275
rect 14685 250 14790 275
rect 17185 250 17290 275
rect 19685 250 19790 275
rect 22185 250 22290 275
rect 24685 250 24790 275
rect 27185 250 27290 275
rect 29685 250 29790 275
rect 32185 250 32290 275
rect 34685 250 34790 275
rect 37185 250 37290 275
rect 39685 250 39790 275
rect 42185 250 42290 275
rect 44685 250 44790 275
rect 47185 250 47290 275
rect -6490 75 -6465 95
rect -4890 75 -4865 95
rect -3290 75 -3265 95
rect -1690 75 -1665 95
rect 740 75 765 95
rect 2340 75 2365 95
rect 3940 75 3965 95
rect 5540 75 5565 95
rect 7970 75 7995 95
rect 9570 75 9595 95
rect 11170 75 11195 95
rect 12770 75 12795 95
rect 15200 75 15225 95
rect 16800 75 16825 95
rect 18400 75 18425 95
rect 20000 75 20025 95
rect 22430 75 22455 95
rect 24030 75 24055 95
rect 25630 75 25655 95
rect 27230 75 27255 95
rect 29660 75 29685 95
rect 31260 75 31285 95
rect 32860 75 32885 95
rect 34460 75 34485 95
rect 36890 75 36915 95
rect 38490 75 38515 95
rect 40090 75 40115 95
rect 41690 75 41715 95
rect 44120 75 44145 95
rect 45720 75 45745 95
rect -10415 15 -9645 35
rect -9615 15 -8845 35
rect 47395 15 48165 35
rect -10415 -295 -9645 -275
rect -9615 -295 -8845 -275
rect 43365 -295 44135 -275
rect 44160 -295 44930 -275
<< metal1 >>
rect -10460 275 48280 315
rect -10460 250 -7815 275
rect -7710 250 -5315 275
rect -5210 250 -2815 275
rect -2710 250 -315 275
rect -210 250 2185 275
rect 2290 250 4685 275
rect 4790 250 7185 275
rect 7290 250 9685 275
rect 9790 250 12185 275
rect 12290 250 14685 275
rect 14790 250 17185 275
rect 17290 250 19685 275
rect 19790 250 22185 275
rect 22290 250 24685 275
rect 24790 250 27185 275
rect 27290 250 29685 275
rect 29790 250 32185 275
rect 32290 250 34685 275
rect 34790 250 37185 275
rect 37290 250 39685 275
rect 39790 250 42185 275
rect 42290 250 44685 275
rect 44790 250 47185 275
rect 47290 250 48280 275
rect -10460 195 48280 250
rect -10460 95 47355 135
rect -10460 75 -6490 95
rect -6465 75 -4890 95
rect -4865 75 -3290 95
rect -3265 75 -1690 95
rect -1665 75 740 95
rect 765 75 2340 95
rect 2365 75 3940 95
rect 3965 75 5540 95
rect 5565 75 7970 95
rect 7995 75 9570 95
rect 9595 75 11170 95
rect 11195 75 12770 95
rect 12795 75 15200 95
rect 15225 75 16800 95
rect 16825 75 18400 95
rect 18425 75 20000 95
rect 20025 75 22430 95
rect 22455 75 24030 95
rect 24055 75 25630 95
rect 25655 75 27230 95
rect 27255 75 29660 95
rect 29685 75 31260 95
rect 31285 75 32860 95
rect 32885 75 34460 95
rect 34485 75 36890 95
rect 36915 75 38490 95
rect 38515 75 40090 95
rect 40115 75 41690 95
rect 41715 75 44120 95
rect 44145 75 45720 95
rect 45745 75 47355 95
rect -10460 65 47355 75
rect -9630 45 -8830 50
rect -10425 35 -8830 45
rect -10425 15 -10415 35
rect -9645 15 -9615 35
rect -8845 15 -8830 35
rect -10425 5 -8830 15
rect 47385 35 48175 45
rect 47385 15 47395 35
rect 48165 15 48175 35
rect 47385 5 48175 15
rect -9630 0 -8830 5
rect -9615 -100 -9590 0
rect 47775 -100 47800 5
rect -10460 -135 47800 -100
rect -9615 -260 -9590 -135
rect -9630 -265 -8830 -260
rect 43745 -265 43770 -135
rect 48215 -265 48280 195
rect -10425 -275 -8830 -265
rect -10425 -295 -10415 -275
rect -9645 -295 -9615 -275
rect -8845 -295 -8830 -275
rect -10425 -305 -8830 -295
rect 43355 -275 48280 -265
rect 43355 -295 43365 -275
rect 44135 -295 44160 -275
rect 44930 -295 48280 -275
rect 43355 -305 48280 -295
rect -9630 -310 -8830 -305
<< labels >>
rlabel locali -3285 -640 -3285 -640 5 V6
port 1 s
rlabel locali -2425 -640 -2425 -640 5 V6i
port 2 s
rlabel locali 3945 -640 3945 -640 5 V5
port 3 s
rlabel locali 4805 -640 4805 -640 5 V5i
port 4 s
rlabel locali 11175 -640 11175 -640 5 V4
port 5 s
rlabel locali 12035 -640 12035 -640 5 V4i
port 6 s
rlabel locali 18405 -640 18405 -640 5 V3
port 7 s
rlabel locali 19265 -640 19265 -640 5 V3i
port 8 s
rlabel locali 25635 -640 25635 -640 5 V2
port 9 s
rlabel locali 26495 -640 26495 -640 5 V2i
port 10 s
rlabel locali 32865 -640 32865 -640 5 V1
port 11 s
rlabel locali 33725 -640 33725 -640 5 V1i
port 12 s
rlabel locali 40095 -640 40095 -640 5 V0
port 13 s
rlabel locali 40955 -640 40955 -640 5 V0i
port 14 s
rlabel locali 48210 -500 48210 -500 3 Idump
port 16 e
rlabel locali 48210 -540 48210 -540 3 Iout
port 17 e
rlabel metal1 -10460 -120 -10460 -120 7 VN
port 18 w
rlabel metal1 -10460 80 -10460 80 7 VP
port 19 w
rlabel locali -10460 195 -10460 195 7 Iin
port 15 w
<< end >>
