* NGSPICE file created from curgen_1.ext - technology: sky130A

X0 a_n1440_n3190# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=96 pd=40 as=48 ps=20 w=12 l=8
X1 a_n3040_n3090# VN VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X2 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X3 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X4 VN VN a_n3040_n3090# VN sky130_fd_pr__nfet_01v8 ad=95.9 pd=40 as=48 ps=20 w=12 l=8
X5 VN a_23200_n100# a_23200_n100# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X6 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X7 a_n3040_n3090# a_n3040_n3090# VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X8 VP Vbp a_n1440_n3190# VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X9 Vbp a_n3040_n3090# VP VP sky130_fd_pr__pfet_01v8 ad=96 pd=40 as=48 ps=20 w=12 l=8
X10 VN a_n1440_n3190# a_n3040_n3090# VN sky130_fd_pr__nfet_01v8 ad=96 pd=40 as=48 ps=20 w=12 l=8
X11 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X12 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X13 a_n3040_n3090# a_n1440_n3190# VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X14 VP Vbp Iin VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X15 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X16 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X17 VP Vbp a_23200_n100# VP sky130_fd_pr__pfet_01v8 ad=96 pd=40 as=48 ps=20 w=12 l=8
X18 VN a_23200_n100# Vbp VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X19 a_23200_n100# a_23200_n100# VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X20 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X21 Vbp VP VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X22 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X23 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=95.9 pd=40 as=48 ps=20 w=12 l=8
X24 Vbp a_23200_n100# VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X25 VN VN Vbp VN sky130_fd_pr__nfet_01v8 ad=90.5 pd=41 as=48 ps=20 w=12 l=8
X26 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X27 a_23200_n100# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X28 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=96 ps=40 w=12 l=8
X29 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X30 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X31 Ires a_n1440_n3190# a_n1440_n3190# VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X32 VP a_n3040_n3090# Vbp VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X33 VP a_n3040_n3090# a_n3040_n3090# VP sky130_fd_pr__pfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X34 a_n1440_n3190# a_n1440_n3190# Ires VN sky130_fd_pr__nfet_01v8 ad=48 pd=20 as=48 ps=20 w=12 l=8
X35 Iin Vbp VP VP sky130_fd_pr__pfet_01v8 ad=96 pd=40 as=48 ps=20 w=12 l=8

