magic
tech sky130A
timestamp 1700264934
<< nwell >>
rect -2460 1640 33780 2525
rect -2460 1600 16060 1640
rect -2460 885 13725 1600
<< nmos >>
rect 16890 805 17690 1405
rect 19320 805 20120 1405
rect 20920 805 21720 1405
rect 22520 805 23320 1405
rect 24120 805 24920 1405
rect 26550 805 27350 1405
rect 28150 805 28950 1405
rect -1600 0 -800 600
rect 0 0 800 600
rect 2430 0 3230 600
rect 4030 0 4830 600
rect 6460 0 7260 600
rect 8060 0 8860 600
rect 10490 0 11290 600
rect 12090 0 12890 600
rect 13690 0 14490 600
rect 15290 0 16090 600
rect 16890 0 17690 600
rect 18490 0 19290 600
rect 20920 0 21720 600
rect 22520 0 23320 600
rect 24950 0 25750 600
rect 26550 0 27350 600
rect 28980 0 29780 600
rect 30580 0 31380 600
<< pmos >>
rect -830 1675 -30 2275
rect 770 1675 1570 2275
rect 3200 1675 4000 2275
rect 4800 1675 5600 2275
rect 7230 1675 8030 2275
rect 8830 1675 9630 2275
rect 11260 1675 12060 2275
rect 12860 1675 13660 2275
rect 14460 1675 15260 2275
rect 16060 1675 16860 2275
rect 17660 1675 18460 2275
rect 19260 1675 20060 2275
rect 21690 1675 22490 2275
rect 23290 1675 24090 2275
rect 25720 1675 26520 2275
rect 27320 1675 28120 2275
rect 29750 1675 30550 2275
rect 31350 1675 32150 2275
rect -830 905 -30 1505
rect 770 905 1570 1505
rect 3200 905 4000 1505
rect 5630 905 6430 1505
rect 7230 905 8030 1505
rect 9660 905 10460 1505
rect 12090 905 12890 1505
<< ndiff >>
rect 16090 1390 16890 1405
rect 16090 820 16105 1390
rect 16875 820 16890 1390
rect 16090 805 16890 820
rect 17690 1390 18490 1405
rect 17690 820 17705 1390
rect 18475 820 18490 1390
rect 17690 805 18490 820
rect 18520 1390 19320 1405
rect 18520 820 18535 1390
rect 19305 820 19320 1390
rect 18520 805 19320 820
rect 20120 1390 20920 1405
rect 20120 820 20135 1390
rect 20905 820 20920 1390
rect 20120 805 20920 820
rect 21720 1390 22520 1405
rect 21720 820 21735 1390
rect 22505 820 22520 1390
rect 21720 805 22520 820
rect 23320 1390 24120 1405
rect 23320 820 23335 1390
rect 24105 820 24120 1390
rect 23320 805 24120 820
rect 24920 1390 25720 1405
rect 24920 820 24935 1390
rect 25705 820 25720 1390
rect 24920 805 25720 820
rect 25750 1390 26550 1405
rect 25750 820 25765 1390
rect 26535 820 26550 1390
rect 25750 805 26550 820
rect 27350 1390 28150 1405
rect 27350 820 27365 1390
rect 28135 820 28150 1390
rect 27350 805 28150 820
rect 28950 1390 29750 1405
rect 28950 820 28965 1390
rect 29735 820 29750 1390
rect 28950 805 29750 820
rect -2400 585 -1600 600
rect -2400 15 -2385 585
rect -1615 15 -1600 585
rect -2400 0 -1600 15
rect -800 585 0 600
rect -800 15 -785 585
rect -15 15 0 585
rect -800 0 0 15
rect 800 585 1600 600
rect 800 15 815 585
rect 1585 15 1600 585
rect 800 0 1600 15
rect 1630 585 2430 600
rect 1630 15 1645 585
rect 2415 15 2430 585
rect 1630 0 2430 15
rect 3230 585 4030 600
rect 3230 15 3245 585
rect 4015 15 4030 585
rect 3230 0 4030 15
rect 4830 585 5630 600
rect 4830 15 4845 585
rect 5615 15 5630 585
rect 4830 0 5630 15
rect 5660 585 6460 600
rect 5660 15 5675 585
rect 6445 15 6460 585
rect 5660 0 6460 15
rect 7260 585 8060 600
rect 7260 15 7275 585
rect 8045 15 8060 585
rect 7260 0 8060 15
rect 8860 585 9660 600
rect 8860 15 8875 585
rect 9645 15 9660 585
rect 8860 0 9660 15
rect 9690 585 10490 600
rect 9690 15 9705 585
rect 10475 15 10490 585
rect 9690 0 10490 15
rect 11290 585 12090 600
rect 11290 15 11305 585
rect 12075 15 12090 585
rect 11290 0 12090 15
rect 12890 585 13690 600
rect 12890 15 12905 585
rect 13675 15 13690 585
rect 12890 0 13690 15
rect 14490 585 15290 600
rect 14490 15 14505 585
rect 15275 15 15290 585
rect 14490 0 15290 15
rect 16090 585 16890 600
rect 16090 15 16105 585
rect 16875 15 16890 585
rect 16090 0 16890 15
rect 17690 585 18490 600
rect 17690 15 17705 585
rect 18475 15 18490 585
rect 17690 0 18490 15
rect 19290 585 20090 600
rect 19290 15 19305 585
rect 20075 15 20090 585
rect 19290 0 20090 15
rect 20120 585 20920 600
rect 20120 15 20135 585
rect 20905 15 20920 585
rect 20120 0 20920 15
rect 21720 585 22520 600
rect 21720 15 21735 585
rect 22505 15 22520 585
rect 21720 0 22520 15
rect 23320 585 24120 600
rect 23320 15 23335 585
rect 24105 15 24120 585
rect 23320 0 24120 15
rect 24150 585 24950 600
rect 24150 15 24165 585
rect 24935 15 24950 585
rect 24150 0 24950 15
rect 25750 585 26550 600
rect 25750 15 25765 585
rect 26535 15 26550 585
rect 25750 0 26550 15
rect 27350 585 28150 600
rect 27350 15 27365 585
rect 28135 15 28150 585
rect 27350 0 28150 15
rect 28180 585 28980 600
rect 28180 15 28195 585
rect 28965 15 28980 585
rect 28180 0 28980 15
rect 29780 585 30580 600
rect 29780 15 29795 585
rect 30565 15 30580 585
rect 29780 0 30580 15
rect 31380 585 32180 600
rect 31380 15 31395 585
rect 32165 15 32180 585
rect 31380 0 32180 15
<< pdiff >>
rect -1630 2260 -830 2275
rect -1630 1690 -1615 2260
rect -845 1690 -830 2260
rect -1630 1675 -830 1690
rect -30 2260 770 2275
rect -30 1690 -15 2260
rect 755 1690 770 2260
rect -30 1675 770 1690
rect 1570 2260 2370 2275
rect 1570 1690 1585 2260
rect 2355 1690 2370 2260
rect 1570 1675 2370 1690
rect 2400 2260 3200 2275
rect 2400 1690 2415 2260
rect 3185 1690 3200 2260
rect 2400 1675 3200 1690
rect 4000 2260 4800 2275
rect 4000 1690 4015 2260
rect 4785 1690 4800 2260
rect 4000 1675 4800 1690
rect 5600 2260 6400 2275
rect 5600 1690 5615 2260
rect 6385 1690 6400 2260
rect 5600 1675 6400 1690
rect 6430 2260 7230 2275
rect 6430 1690 6445 2260
rect 7215 1690 7230 2260
rect 6430 1675 7230 1690
rect 8030 2260 8830 2275
rect 8030 1690 8045 2260
rect 8815 1690 8830 2260
rect 8030 1675 8830 1690
rect 9630 2260 10430 2275
rect 9630 1690 9645 2260
rect 10415 1690 10430 2260
rect 9630 1675 10430 1690
rect 10460 2260 11260 2275
rect 10460 1690 10475 2260
rect 11245 1690 11260 2260
rect 10460 1675 11260 1690
rect 12060 2260 12860 2275
rect 12060 1690 12075 2260
rect 12845 1690 12860 2260
rect 12060 1675 12860 1690
rect 13660 2260 14460 2275
rect 13660 1690 13675 2260
rect 14445 1690 14460 2260
rect 13660 1675 14460 1690
rect 15260 2260 16060 2275
rect 15260 1690 15275 2260
rect 16045 1690 16060 2260
rect 15260 1675 16060 1690
rect 16860 2260 17660 2275
rect 16860 1690 16875 2260
rect 17645 1690 17660 2260
rect 16860 1675 17660 1690
rect 18460 2260 19260 2275
rect 18460 1690 18475 2260
rect 19245 1690 19260 2260
rect 18460 1675 19260 1690
rect 20060 2260 20860 2275
rect 20060 1690 20075 2260
rect 20845 1690 20860 2260
rect 20060 1675 20860 1690
rect 20890 2260 21690 2275
rect 20890 1690 20905 2260
rect 21675 1690 21690 2260
rect 20890 1675 21690 1690
rect 22490 2260 23290 2275
rect 22490 1690 22505 2260
rect 23275 1690 23290 2260
rect 22490 1675 23290 1690
rect 24090 2260 24890 2275
rect 24090 1690 24105 2260
rect 24875 1690 24890 2260
rect 24090 1675 24890 1690
rect 24920 2260 25720 2275
rect 24920 1690 24935 2260
rect 25705 1690 25720 2260
rect 24920 1675 25720 1690
rect 26520 2260 27320 2275
rect 26520 1690 26535 2260
rect 27305 1690 27320 2260
rect 26520 1675 27320 1690
rect 28120 2260 28920 2275
rect 28120 1690 28135 2260
rect 28905 1690 28920 2260
rect 28120 1675 28920 1690
rect 28950 2260 29750 2275
rect 28950 1690 28965 2260
rect 29735 1690 29750 2260
rect 28950 1675 29750 1690
rect 30550 2260 31350 2275
rect 30550 1690 30565 2260
rect 31335 1690 31350 2260
rect 30550 1675 31350 1690
rect 32150 2260 32950 2275
rect 32150 1690 32165 2260
rect 32935 1690 32950 2260
rect 32150 1675 32950 1690
rect -1630 1490 -830 1505
rect -1630 920 -1615 1490
rect -845 920 -830 1490
rect -1630 905 -830 920
rect -30 1490 770 1505
rect -30 920 -15 1490
rect 755 920 770 1490
rect -30 905 770 920
rect 1570 1490 2370 1505
rect 1570 920 1585 1490
rect 2355 920 2370 1490
rect 1570 905 2370 920
rect 2400 1490 3200 1505
rect 2400 920 2415 1490
rect 3185 920 3200 1490
rect 2400 905 3200 920
rect 4000 1490 4800 1505
rect 4000 920 4015 1490
rect 4785 920 4800 1490
rect 4000 905 4800 920
rect 4830 1490 5630 1505
rect 4830 920 4845 1490
rect 5615 920 5630 1490
rect 4830 905 5630 920
rect 6430 1490 7230 1505
rect 6430 920 6445 1490
rect 7215 920 7230 1490
rect 6430 905 7230 920
rect 8030 1490 8830 1505
rect 8030 920 8045 1490
rect 8815 920 8830 1490
rect 8030 905 8830 920
rect 8860 1490 9660 1505
rect 8860 920 8875 1490
rect 9645 920 9660 1490
rect 8860 905 9660 920
rect 10460 1490 11260 1505
rect 10460 920 10475 1490
rect 11245 920 11260 1490
rect 10460 905 11260 920
rect 11290 1490 12090 1505
rect 11290 920 11305 1490
rect 12075 920 12090 1490
rect 11290 905 12090 920
rect 12890 1490 13690 1505
rect 12890 920 12905 1490
rect 13675 920 13690 1490
rect 12890 905 13690 920
<< ndiffc >>
rect 16105 820 16875 1390
rect 17705 820 18475 1390
rect 18535 820 19305 1390
rect 20135 820 20905 1390
rect 21735 820 22505 1390
rect 23335 820 24105 1390
rect 24935 820 25705 1390
rect 25765 820 26535 1390
rect 27365 820 28135 1390
rect 28965 820 29735 1390
rect -2385 15 -1615 585
rect -785 15 -15 585
rect 815 15 1585 585
rect 1645 15 2415 585
rect 3245 15 4015 585
rect 4845 15 5615 585
rect 5675 15 6445 585
rect 7275 15 8045 585
rect 8875 15 9645 585
rect 9705 15 10475 585
rect 11305 15 12075 585
rect 12905 15 13675 585
rect 14505 15 15275 585
rect 16105 15 16875 585
rect 17705 15 18475 585
rect 19305 15 20075 585
rect 20135 15 20905 585
rect 21735 15 22505 585
rect 23335 15 24105 585
rect 24165 15 24935 585
rect 25765 15 26535 585
rect 27365 15 28135 585
rect 28195 15 28965 585
rect 29795 15 30565 585
rect 31395 15 32165 585
<< pdiffc >>
rect -1615 1690 -845 2260
rect -15 1690 755 2260
rect 1585 1690 2355 2260
rect 2415 1690 3185 2260
rect 4015 1690 4785 2260
rect 5615 1690 6385 2260
rect 6445 1690 7215 2260
rect 8045 1690 8815 2260
rect 9645 1690 10415 2260
rect 10475 1690 11245 2260
rect 12075 1690 12845 2260
rect 13675 1690 14445 2260
rect 15275 1690 16045 2260
rect 16875 1690 17645 2260
rect 18475 1690 19245 2260
rect 20075 1690 20845 2260
rect 20905 1690 21675 2260
rect 22505 1690 23275 2260
rect 24105 1690 24875 2260
rect 24935 1690 25705 2260
rect 26535 1690 27305 2260
rect 28135 1690 28905 2260
rect 28965 1690 29735 2260
rect 30565 1690 31335 2260
rect 32165 1690 32935 2260
rect -1615 920 -845 1490
rect -15 920 755 1490
rect 1585 920 2355 1490
rect 2415 920 3185 1490
rect 4015 920 4785 1490
rect 4845 920 5615 1490
rect 6445 920 7215 1490
rect 8045 920 8815 1490
rect 8875 920 9645 1490
rect 10475 920 11245 1490
rect 11305 920 12075 1490
rect 12905 920 13675 1490
<< psubdiff >>
rect 29750 1390 30550 1405
rect 29750 820 29765 1390
rect 30535 820 30550 1390
rect 29750 805 30550 820
rect -3200 585 -2400 600
rect -3200 15 -3185 585
rect -2415 15 -2400 585
rect -3200 0 -2400 15
rect 32180 585 32980 600
rect 32180 15 32195 585
rect 32965 15 32980 585
rect 32180 0 32980 15
<< nsubdiff >>
rect -2430 2260 -1630 2275
rect -2430 1690 -2415 2260
rect -1645 1690 -1630 2260
rect -2430 1675 -1630 1690
rect 32950 2260 33750 2275
rect 32950 1690 32965 2260
rect 33735 1690 33750 2260
rect 32950 1675 33750 1690
rect -2430 1490 -1630 1505
rect -2430 920 -2415 1490
rect -1645 920 -1630 1490
rect -2430 905 -1630 920
<< psubdiffcont >>
rect 29765 820 30535 1390
rect -3185 15 -2415 585
rect 32195 15 32965 585
<< nsubdiffcont >>
rect -2415 1690 -1645 2260
rect 32965 1690 33735 2260
rect -2415 920 -1645 1490
<< poly >>
rect 7455 2465 7500 2475
rect 7455 2445 7465 2465
rect 7490 2445 7500 2465
rect 7455 2440 7500 2445
rect 11545 2465 11590 2475
rect 11545 2445 11555 2465
rect 11580 2445 11590 2465
rect 11545 2440 11590 2445
rect 19730 2465 19775 2470
rect 19730 2445 19740 2465
rect 19765 2445 19775 2465
rect 19730 2440 19775 2445
rect 23820 2465 23865 2470
rect 23820 2445 23830 2465
rect 23855 2445 23865 2465
rect 23820 2440 23865 2445
rect -810 2340 -765 2350
rect -810 2320 -800 2340
rect -775 2320 -765 2340
rect -810 2315 -765 2320
rect 790 2340 835 2350
rect 790 2320 800 2340
rect 825 2320 835 2340
rect 790 2315 835 2320
rect 3220 2340 3265 2350
rect 3220 2320 3230 2340
rect 3255 2320 3265 2340
rect 3220 2315 3265 2320
rect 4820 2340 4865 2350
rect 4820 2320 4830 2340
rect 4855 2320 4865 2340
rect 4820 2315 4865 2320
rect 6605 2340 6650 2350
rect 6605 2320 6615 2340
rect 6640 2330 6650 2340
rect 6755 2340 6800 2350
rect 6755 2330 6765 2340
rect 6640 2320 6765 2330
rect 6790 2320 6800 2340
rect 6605 2315 6800 2320
rect -805 2290 -790 2315
rect 795 2290 810 2315
rect 3225 2290 3240 2315
rect 4825 2290 4840 2315
rect 7470 2290 7485 2440
rect 8850 2340 8895 2350
rect 8850 2320 8860 2340
rect 8885 2320 8895 2340
rect 8850 2315 8895 2320
rect 10575 2340 10620 2350
rect 10575 2320 10585 2340
rect 10610 2330 10620 2340
rect 10725 2340 10770 2350
rect 10725 2330 10735 2340
rect 10610 2320 10735 2330
rect 10760 2320 10770 2340
rect 10575 2315 10770 2320
rect 8855 2290 8870 2315
rect 11560 2290 11575 2440
rect 12880 2340 12925 2350
rect 12880 2320 12890 2340
rect 12915 2320 12925 2340
rect 12880 2315 12925 2320
rect 14480 2340 14525 2350
rect 14480 2320 14490 2340
rect 14515 2320 14525 2340
rect 14480 2315 14525 2320
rect 16795 2340 16840 2350
rect 16795 2320 16805 2340
rect 16830 2320 16840 2340
rect 16795 2315 16840 2320
rect 18395 2340 18440 2350
rect 18395 2320 18405 2340
rect 18430 2320 18440 2340
rect 18395 2315 18440 2320
rect 12885 2290 12905 2315
rect 14485 2290 14505 2315
rect 16815 2290 16835 2315
rect 18415 2290 18435 2315
rect 19745 2290 19760 2440
rect 20550 2340 20595 2350
rect 20550 2320 20560 2340
rect 20585 2330 20595 2340
rect 20700 2340 20745 2350
rect 20700 2330 20710 2340
rect 20585 2320 20710 2330
rect 20735 2320 20745 2340
rect 20550 2315 20745 2320
rect 22425 2340 22470 2350
rect 22425 2320 22435 2340
rect 22460 2320 22470 2340
rect 22425 2315 22470 2320
rect 22450 2290 22465 2315
rect 23835 2290 23850 2440
rect 33715 2400 33760 2410
rect 33715 2380 33725 2400
rect 33750 2390 33760 2400
rect 33885 2400 33930 2410
rect 33885 2390 33895 2400
rect 33750 2380 33895 2390
rect 33920 2380 33930 2400
rect 33715 2375 33930 2380
rect 24520 2340 24565 2350
rect 24520 2320 24530 2340
rect 24555 2330 24565 2340
rect 24670 2340 24715 2350
rect 24670 2330 24680 2340
rect 24555 2320 24680 2330
rect 24705 2320 24715 2340
rect 24520 2315 24715 2320
rect 26455 2340 26500 2350
rect 26455 2320 26465 2340
rect 26490 2320 26500 2340
rect 26455 2315 26500 2320
rect 28055 2340 28100 2350
rect 28055 2320 28065 2340
rect 28090 2320 28100 2340
rect 28055 2315 28100 2320
rect 30485 2340 30530 2350
rect 30485 2320 30495 2340
rect 30520 2320 30530 2340
rect 30485 2315 30530 2320
rect 32085 2340 32130 2350
rect 32085 2320 32095 2340
rect 32120 2320 32130 2340
rect 32085 2315 32130 2320
rect 26480 2290 26495 2315
rect 28080 2290 28095 2315
rect 30510 2290 30525 2315
rect 32110 2290 32125 2315
rect -830 2275 -30 2290
rect 770 2275 1570 2290
rect 3200 2275 4000 2290
rect 4800 2275 5600 2290
rect 7230 2275 8030 2290
rect 8830 2275 9630 2290
rect 11260 2275 12060 2290
rect 12860 2275 13660 2290
rect 14460 2275 15260 2290
rect 16060 2275 16860 2290
rect 17660 2275 18460 2290
rect 19260 2275 20060 2290
rect 21690 2275 22490 2290
rect 23290 2275 24090 2290
rect 25720 2275 26520 2290
rect 27320 2275 28120 2290
rect 29750 2275 30550 2290
rect 31350 2275 32150 2290
rect -830 1660 -30 1675
rect 770 1660 1570 1675
rect 3200 1660 4000 1675
rect 4800 1660 5600 1675
rect 7230 1660 8030 1675
rect 8830 1660 9630 1675
rect 11260 1660 12060 1675
rect 12860 1660 13660 1675
rect 14460 1660 15260 1675
rect 16060 1660 16860 1675
rect 17660 1660 18460 1675
rect 19260 1660 20060 1675
rect 21690 1660 22490 1675
rect 23290 1660 24090 1675
rect 25720 1660 26520 1675
rect 27320 1660 28120 1675
rect 29750 1660 30550 1675
rect 31350 1660 32150 1675
rect -805 1570 -760 1580
rect -805 1550 -795 1570
rect -770 1550 -760 1570
rect -805 1545 -760 1550
rect 1525 1570 1570 1580
rect 1525 1550 1535 1570
rect 1560 1550 1570 1570
rect 1525 1545 1570 1550
rect 2850 1570 2895 1580
rect 2850 1550 2860 1570
rect 2885 1560 2895 1570
rect 3000 1570 3045 1580
rect 3000 1560 3010 1570
rect 2885 1550 3010 1560
rect 3035 1550 3045 1570
rect 2850 1545 3045 1550
rect 3955 1570 4000 1580
rect 3955 1550 3965 1570
rect 3990 1550 4000 1570
rect 3955 1545 4000 1550
rect 4955 1570 5000 1580
rect 4955 1550 4965 1570
rect 4990 1560 5000 1570
rect 5105 1570 5150 1580
rect 5105 1560 5115 1570
rect 4990 1550 5115 1560
rect 5140 1550 5150 1570
rect 4955 1545 5150 1550
rect 6385 1570 6430 1580
rect 6385 1550 6395 1570
rect 6420 1550 6430 1570
rect 6385 1545 6430 1550
rect -800 1520 -785 1545
rect 1555 1520 1570 1545
rect 3985 1520 4000 1545
rect 6415 1520 6430 1545
rect -830 1505 -30 1520
rect 770 1505 1570 1520
rect 3200 1505 4000 1520
rect 5630 1505 6430 1520
rect 7230 1570 7275 1580
rect 7230 1550 7240 1570
rect 7265 1550 7275 1570
rect 7230 1545 7275 1550
rect 8510 1570 8555 1580
rect 8510 1550 8520 1570
rect 8545 1560 8555 1570
rect 8660 1570 8705 1580
rect 8660 1560 8670 1570
rect 8545 1550 8670 1560
rect 8695 1550 8705 1570
rect 8510 1545 8705 1550
rect 9660 1570 9705 1580
rect 9660 1550 9670 1570
rect 9695 1550 9705 1570
rect 9660 1545 9705 1550
rect 10615 1570 10660 1580
rect 10615 1550 10625 1570
rect 10650 1560 10660 1570
rect 10765 1570 10810 1580
rect 10765 1560 10775 1570
rect 10650 1550 10775 1560
rect 10800 1550 10810 1570
rect 10615 1545 10810 1550
rect 12090 1570 12135 1580
rect 12090 1550 12100 1570
rect 12125 1550 12135 1570
rect 12090 1545 12135 1550
rect 7230 1520 7245 1545
rect 9660 1520 9675 1545
rect 12090 1520 12105 1545
rect 7230 1505 8030 1520
rect 9660 1505 10460 1520
rect 12090 1505 12890 1520
rect 21625 1485 21875 1495
rect 21625 1465 21635 1485
rect 21660 1480 21840 1485
rect 21660 1465 21670 1480
rect 21625 1460 21670 1465
rect 21830 1465 21840 1480
rect 21865 1465 21875 1485
rect 21830 1460 21875 1465
rect 16890 1405 17690 1420
rect 19320 1405 20120 1420
rect 20920 1405 21720 1420
rect 22520 1405 23320 1420
rect 24120 1405 24920 1420
rect 26550 1405 27350 1420
rect 28150 1405 28950 1420
rect -830 890 -30 905
rect 770 890 1570 905
rect 3200 890 4000 905
rect 5630 890 6430 905
rect 7230 890 8030 905
rect 9660 890 10460 905
rect 12090 890 12890 905
rect 6745 845 6790 855
rect 6745 825 6755 845
rect 6780 835 6790 845
rect 6930 845 6975 855
rect 6930 835 6940 845
rect 6780 825 6940 835
rect 6965 825 6975 845
rect 6745 820 6975 825
rect 16890 790 17690 805
rect 19320 790 20120 805
rect 20920 790 21720 805
rect 22520 790 23320 805
rect 24120 790 24920 805
rect 26550 790 27350 805
rect 28150 790 28950 805
rect 6745 780 6790 790
rect 6745 760 6755 780
rect 6780 770 6790 780
rect 6930 780 6975 790
rect 6930 770 6940 780
rect 6780 760 6940 770
rect 6965 760 6975 780
rect 6745 755 6975 760
rect 9050 780 9095 790
rect 9050 760 9060 780
rect 9085 770 9095 780
rect 9215 780 9260 790
rect 9215 770 9225 780
rect 9085 760 9225 770
rect 9250 760 9260 780
rect 9050 755 9260 760
rect 16890 785 16935 790
rect 16890 765 16900 785
rect 16925 765 16935 785
rect 16890 755 16935 765
rect 19320 785 19365 790
rect 19320 765 19330 785
rect 19355 765 19365 785
rect 19320 755 19365 765
rect 20920 785 20965 790
rect 20920 765 20930 785
rect 20955 765 20965 785
rect 20920 755 20965 765
rect 23275 785 23320 790
rect 23275 765 23285 785
rect 23310 765 23320 785
rect 23275 755 23320 765
rect 24875 785 24920 790
rect 24875 765 24885 785
rect 24910 765 24920 785
rect 24875 755 24920 765
rect 27305 785 27350 790
rect 27305 765 27315 785
rect 27340 765 27350 785
rect 27305 755 27350 765
rect 28880 785 28925 790
rect 28880 765 28890 785
rect 28915 765 28925 785
rect 28880 755 28925 765
rect 6460 720 6505 730
rect 6460 700 6470 720
rect 6495 700 6505 720
rect 6460 695 6505 700
rect 6745 720 6790 730
rect 6745 700 6755 720
rect 6780 710 6790 720
rect 6930 720 6975 730
rect 6930 710 6940 720
rect 6780 700 6940 710
rect 6965 700 6975 720
rect 6745 695 6975 700
rect 10490 720 10535 730
rect 10490 700 10500 720
rect 10525 700 10535 720
rect 10490 695 10535 700
rect 19245 720 19290 730
rect 19245 700 19255 720
rect 19280 700 19290 720
rect 19245 695 19290 700
rect 23275 720 23320 730
rect 23275 700 23285 720
rect 23310 700 23320 720
rect 23275 695 23320 700
rect 0 665 45 675
rect 0 645 10 665
rect 35 645 45 665
rect 0 640 45 645
rect 2430 665 2475 675
rect 2430 645 2440 665
rect 2465 645 2475 665
rect 2430 640 2475 645
rect 4030 665 4075 675
rect 4030 645 4040 665
rect 4065 645 4075 665
rect 4030 640 4075 645
rect 5590 665 5635 675
rect 5590 645 5600 665
rect 5625 655 5635 665
rect 5740 665 5785 675
rect 5740 655 5750 665
rect 5625 645 5750 655
rect 5775 645 5785 665
rect 5590 640 5785 645
rect 0 615 15 640
rect 2430 615 2445 640
rect 4030 615 4045 640
rect 6460 615 6475 695
rect 8060 665 8105 675
rect 8060 645 8070 665
rect 8095 645 8105 665
rect 8060 640 8105 645
rect 9620 665 9665 675
rect 9620 645 9630 665
rect 9655 655 9665 665
rect 9770 665 9815 675
rect 9770 655 9780 665
rect 9655 645 9780 655
rect 9805 645 9815 665
rect 9620 640 9815 645
rect 8060 615 8075 640
rect 10490 615 10505 695
rect 12090 665 12135 675
rect 12090 645 12100 665
rect 12125 645 12135 665
rect 12090 640 12135 645
rect 13690 665 13735 675
rect 13690 645 13700 665
rect 13725 645 13735 665
rect 13690 640 13735 645
rect 16045 665 16090 675
rect 16045 645 16055 665
rect 16080 645 16090 665
rect 16045 640 16090 645
rect 17645 665 17690 675
rect 17645 645 17655 665
rect 17680 645 17690 665
rect 17645 640 17690 645
rect 12090 615 12105 640
rect 13690 615 13705 640
rect 16075 615 16090 640
rect 17675 615 17690 640
rect 19275 615 19290 695
rect 19965 665 20010 675
rect 19965 645 19975 665
rect 20000 655 20010 665
rect 20115 665 20160 675
rect 20115 655 20125 665
rect 20000 645 20125 655
rect 20150 645 20160 665
rect 19965 640 20160 645
rect 21675 665 21720 675
rect 21675 645 21685 665
rect 21710 645 21720 665
rect 21675 640 21720 645
rect 21705 615 21720 640
rect 23305 615 23320 695
rect 23995 665 24040 675
rect 23995 645 24005 665
rect 24030 655 24040 665
rect 24145 665 24190 675
rect 24145 655 24155 665
rect 24030 645 24155 655
rect 24180 645 24190 665
rect 23995 640 24190 645
rect 25705 665 25750 675
rect 25705 645 25715 665
rect 25740 645 25750 665
rect 25705 640 25750 645
rect 27305 665 27350 675
rect 27305 645 27315 665
rect 27340 645 27350 665
rect 27305 640 27350 645
rect 29735 665 29780 675
rect 29735 645 29745 665
rect 29770 645 29780 665
rect 29735 640 29780 645
rect 25735 615 25750 640
rect 27335 615 27350 640
rect 29765 615 29780 640
rect -1600 600 -800 615
rect 0 600 800 615
rect 2430 600 3230 615
rect 4030 600 4830 615
rect 6460 600 7260 615
rect 8060 600 8860 615
rect 10490 600 11290 615
rect 12090 600 12890 615
rect 13690 600 14490 615
rect 15290 600 16090 615
rect 16890 600 17690 615
rect 18490 600 19290 615
rect 20920 600 21720 615
rect 22520 600 23320 615
rect 24950 600 25750 615
rect 26550 600 27350 615
rect 28980 600 29780 615
rect 30580 600 31380 615
rect -1600 -15 -800 0
rect 0 -15 800 0
rect 2430 -15 3230 0
rect 4030 -15 4830 0
rect 6460 -15 7260 0
rect 8060 -15 8860 0
rect 10490 -15 11290 0
rect 12090 -15 12890 0
rect 13690 -15 14490 0
rect 15290 -15 16090 0
rect 16890 -15 17690 0
rect 18490 -15 19290 0
rect 20920 -15 21720 0
rect 22520 -15 23320 0
rect 24950 -15 25750 0
rect 26550 -15 27350 0
rect 28980 -15 29780 0
rect 30580 -15 31380 0
rect -1600 -20 -1555 -15
rect -1600 -40 -1590 -20
rect -1565 -40 -1555 -20
rect -1600 -50 -1555 -40
rect 31335 -20 31380 -15
rect 31335 -40 31345 -20
rect 31370 -40 31380 -20
rect 31335 -50 31380 -40
<< polycont >>
rect 7465 2445 7490 2465
rect 11555 2445 11580 2465
rect 19740 2445 19765 2465
rect 23830 2445 23855 2465
rect -800 2320 -775 2340
rect 800 2320 825 2340
rect 3230 2320 3255 2340
rect 4830 2320 4855 2340
rect 6615 2320 6640 2340
rect 6765 2320 6790 2340
rect 8860 2320 8885 2340
rect 10585 2320 10610 2340
rect 10735 2320 10760 2340
rect 12890 2320 12915 2340
rect 14490 2320 14515 2340
rect 16805 2320 16830 2340
rect 18405 2320 18430 2340
rect 20560 2320 20585 2340
rect 20710 2320 20735 2340
rect 22435 2320 22460 2340
rect 33725 2380 33750 2400
rect 33895 2380 33920 2400
rect 24530 2320 24555 2340
rect 24680 2320 24705 2340
rect 26465 2320 26490 2340
rect 28065 2320 28090 2340
rect 30495 2320 30520 2340
rect 32095 2320 32120 2340
rect -795 1550 -770 1570
rect 1535 1550 1560 1570
rect 2860 1550 2885 1570
rect 3010 1550 3035 1570
rect 3965 1550 3990 1570
rect 4965 1550 4990 1570
rect 5115 1550 5140 1570
rect 6395 1550 6420 1570
rect 7240 1550 7265 1570
rect 8520 1550 8545 1570
rect 8670 1550 8695 1570
rect 9670 1550 9695 1570
rect 10625 1550 10650 1570
rect 10775 1550 10800 1570
rect 12100 1550 12125 1570
rect 21635 1465 21660 1485
rect 21840 1465 21865 1485
rect 6755 825 6780 845
rect 6940 825 6965 845
rect 6755 760 6780 780
rect 6940 760 6965 780
rect 9060 760 9085 780
rect 9225 760 9250 780
rect 16900 765 16925 785
rect 19330 765 19355 785
rect 20930 765 20955 785
rect 23285 765 23310 785
rect 24885 765 24910 785
rect 27315 765 27340 785
rect 28890 765 28915 785
rect 6470 700 6495 720
rect 6755 700 6780 720
rect 6940 700 6965 720
rect 10500 700 10525 720
rect 19255 700 19280 720
rect 23285 700 23310 720
rect 10 645 35 665
rect 2440 645 2465 665
rect 4040 645 4065 665
rect 5600 645 5625 665
rect 5750 645 5775 665
rect 8070 645 8095 665
rect 9630 645 9655 665
rect 9780 645 9805 665
rect 12100 645 12125 665
rect 13700 645 13725 665
rect 16055 645 16080 665
rect 17655 645 17680 665
rect 19975 645 20000 665
rect 20125 645 20150 665
rect 21685 645 21710 665
rect 24005 645 24030 665
rect 24155 645 24180 665
rect 25715 645 25740 665
rect 27315 645 27340 665
rect 29745 645 29770 665
rect -1590 -40 -1565 -20
rect 31345 -40 31370 -20
<< locali >>
rect 7455 2465 7500 2475
rect 7455 2460 7465 2465
rect 6690 2445 7465 2460
rect 7490 2460 7500 2465
rect 11545 2465 11590 2475
rect 11545 2460 11555 2465
rect 7490 2445 11555 2460
rect 11580 2460 11590 2465
rect 19730 2465 19775 2470
rect 19730 2460 19740 2465
rect 11580 2445 19740 2460
rect 19765 2460 19775 2465
rect 23820 2465 23865 2470
rect 23820 2460 23830 2465
rect 19765 2445 23830 2460
rect 23855 2460 23865 2465
rect 23855 2445 33945 2460
rect 6690 2440 33945 2445
rect -810 2340 -765 2350
rect -810 2335 -800 2340
rect -855 2320 -800 2335
rect -775 2320 -765 2340
rect -855 2315 -765 2320
rect 790 2340 835 2350
rect 790 2320 800 2340
rect 825 2335 835 2340
rect 3220 2340 3265 2350
rect 3220 2335 3230 2340
rect 825 2320 3230 2335
rect 3255 2335 3265 2340
rect 4820 2340 4865 2350
rect 4820 2335 4830 2340
rect 3255 2320 4830 2335
rect 4855 2335 4865 2340
rect 6605 2340 6650 2350
rect 6605 2335 6615 2340
rect 4855 2320 6615 2335
rect 6640 2320 6650 2340
rect 790 2315 6650 2320
rect -855 2270 -835 2315
rect 5605 2270 5625 2315
rect 6690 2270 6710 2440
rect 6755 2340 6800 2350
rect 6755 2320 6765 2340
rect 6790 2335 6800 2340
rect 8850 2340 8895 2350
rect 8850 2335 8860 2340
rect 6790 2320 8860 2335
rect 8885 2335 8895 2340
rect 10575 2340 10620 2350
rect 10575 2335 10585 2340
rect 8885 2320 10585 2335
rect 10610 2320 10620 2340
rect 6755 2315 10620 2320
rect 9635 2270 9655 2315
rect 10660 2270 10680 2440
rect 10725 2340 10770 2350
rect 10725 2320 10735 2340
rect 10760 2335 10770 2340
rect 12880 2340 12925 2350
rect 12880 2335 12890 2340
rect 10760 2320 12890 2335
rect 12915 2335 12925 2340
rect 14480 2340 14525 2350
rect 14480 2335 14490 2340
rect 12915 2320 14490 2335
rect 14515 2335 14525 2340
rect 16795 2340 16840 2350
rect 16795 2335 16805 2340
rect 14515 2320 16805 2335
rect 16830 2335 16840 2340
rect 18395 2340 18440 2350
rect 18395 2335 18405 2340
rect 16830 2320 18405 2335
rect 18430 2335 18440 2340
rect 20550 2340 20595 2350
rect 20550 2335 20560 2340
rect 18430 2320 20560 2335
rect 20585 2320 20595 2340
rect 10725 2315 20595 2320
rect 13665 2270 13685 2315
rect 17635 2270 17655 2315
rect 20640 2270 20660 2440
rect 20700 2340 20745 2350
rect 20700 2320 20710 2340
rect 20735 2335 20745 2340
rect 22425 2340 22470 2350
rect 22425 2335 22435 2340
rect 20735 2320 22435 2335
rect 22460 2335 22470 2340
rect 24520 2340 24565 2350
rect 24520 2335 24530 2340
rect 22460 2320 24530 2335
rect 24555 2320 24565 2340
rect 20700 2315 24565 2320
rect 21665 2270 21685 2315
rect 24610 2270 24630 2440
rect 33715 2400 33760 2410
rect 33715 2395 33725 2400
rect 30510 2380 33725 2395
rect 33750 2380 33760 2400
rect 30510 2375 33760 2380
rect 30510 2350 30530 2375
rect 24670 2340 24715 2350
rect 24670 2320 24680 2340
rect 24705 2335 24715 2340
rect 26455 2340 26500 2350
rect 26455 2335 26465 2340
rect 24705 2320 26465 2335
rect 26490 2335 26500 2340
rect 28055 2340 28100 2350
rect 28055 2335 28065 2340
rect 26490 2320 28065 2335
rect 28090 2335 28100 2340
rect 30485 2340 30530 2350
rect 30485 2335 30495 2340
rect 28090 2320 30495 2335
rect 30520 2320 30530 2340
rect 24670 2315 30530 2320
rect 32085 2340 32130 2350
rect 32085 2320 32095 2340
rect 32120 2335 32130 2340
rect 33740 2335 33760 2375
rect 32120 2320 32175 2335
rect 32085 2315 32175 2320
rect 33740 2315 33815 2335
rect 25695 2270 25715 2315
rect 32155 2270 32175 2315
rect -2425 2260 -835 2270
rect -2425 1690 -2415 2260
rect -1645 1690 -1615 2260
rect -845 1690 -835 2260
rect -2425 1680 -835 1690
rect -25 2260 765 2270
rect -25 1690 -15 2260
rect 755 1690 765 2260
rect -25 1680 765 1690
rect 1575 2260 2365 2270
rect 1575 1690 1585 2260
rect 2355 1690 2365 2260
rect 1575 1680 2365 1690
rect 2405 2260 3195 2270
rect 2405 1690 2415 2260
rect 3185 1690 3195 2260
rect 2405 1680 3195 1690
rect 4005 2260 4795 2270
rect 4005 1690 4015 2260
rect 4785 1690 4795 2260
rect 4005 1680 4795 1690
rect 5605 2260 6395 2270
rect 5605 1690 5615 2260
rect 6385 1690 6395 2260
rect 5605 1680 6395 1690
rect 6435 2260 7225 2270
rect 6435 1690 6445 2260
rect 7215 1690 7225 2260
rect 6435 1680 7225 1690
rect 8035 2260 8825 2270
rect 8035 1690 8045 2260
rect 8815 1690 8825 2260
rect 8035 1680 8825 1690
rect 9635 2260 10425 2270
rect 9635 1690 9645 2260
rect 10415 1690 10425 2260
rect 9635 1680 10425 1690
rect 10465 2260 11255 2270
rect 10465 1690 10475 2260
rect 11245 1690 11255 2260
rect 10465 1680 11255 1690
rect 12065 2260 12855 2270
rect 12065 1690 12075 2260
rect 12845 1690 12855 2260
rect 12065 1680 12855 1690
rect 13665 2260 14455 2270
rect 13665 1690 13675 2260
rect 14445 1690 14455 2260
rect 13665 1680 14455 1690
rect 15265 2260 16055 2270
rect 15265 1690 15275 2260
rect 16045 1690 16055 2260
rect 15265 1680 16055 1690
rect 16865 2260 17655 2270
rect 16865 1690 16875 2260
rect 17645 1690 17655 2260
rect 16865 1680 17655 1690
rect 18465 2260 19255 2270
rect 18465 1690 18475 2260
rect 19245 1690 19255 2260
rect 18465 1680 19255 1690
rect 20065 2260 20855 2270
rect 20065 1690 20075 2260
rect 20845 1690 20855 2260
rect 20065 1680 20855 1690
rect 20895 2260 21685 2270
rect 20895 1690 20905 2260
rect 21675 1690 21685 2260
rect 20895 1680 21685 1690
rect 22495 2260 23285 2270
rect 22495 1690 22505 2260
rect 23275 1690 23285 2260
rect 22495 1680 23285 1690
rect 24095 2260 24885 2270
rect 24095 1690 24105 2260
rect 24875 1690 24885 2260
rect 24095 1680 24885 1690
rect 24925 2260 25715 2270
rect 24925 1690 24935 2260
rect 25705 1690 25715 2260
rect 24925 1680 25715 1690
rect 26525 2260 27315 2270
rect 26525 1690 26535 2260
rect 27305 1690 27315 2260
rect 26525 1680 27315 1690
rect 28125 2260 28915 2270
rect 28125 1690 28135 2260
rect 28905 1690 28915 2260
rect 28125 1680 28915 1690
rect 28955 2260 29745 2270
rect 28955 1690 28965 2260
rect 29735 1690 29745 2260
rect 28955 1680 29745 1690
rect 30555 2260 31345 2270
rect 30555 1690 30565 2260
rect 31335 1690 31345 2260
rect 30555 1680 31345 1690
rect 32155 2260 33745 2270
rect 32155 1690 32165 2260
rect 32935 1690 32965 2260
rect 33735 1690 33745 2260
rect 32155 1680 33745 1690
rect 2345 1660 2365 1680
rect 4775 1660 4795 1680
rect 8805 1660 8825 1680
rect 12380 1660 12400 1680
rect 15670 1660 15690 1680
rect 18920 1660 18940 1680
rect 22495 1660 22515 1680
rect 26525 1660 26545 1680
rect 28955 1660 28975 1680
rect 2345 1640 28975 1660
rect -3230 1605 -685 1625
rect -705 1580 -685 1605
rect -805 1570 -760 1580
rect -805 1550 -795 1570
rect -770 1550 -760 1570
rect -705 1570 1570 1580
rect -705 1560 1535 1570
rect -805 1545 -760 1550
rect 1525 1550 1535 1560
rect 1560 1565 1570 1570
rect 2850 1570 2895 1580
rect 2850 1565 2860 1570
rect 1560 1550 2860 1565
rect 2885 1550 2895 1570
rect 3000 1570 3045 1580
rect 1525 1545 2895 1550
rect -855 1525 -785 1545
rect -855 1500 -835 1525
rect 745 1500 765 1505
rect 2940 1500 2960 1560
rect 3000 1550 3010 1570
rect 3035 1565 3045 1570
rect 3955 1570 4000 1580
rect 3955 1565 3965 1570
rect 3035 1550 3965 1565
rect 3990 1565 4000 1570
rect 4955 1570 5000 1580
rect 4955 1565 4965 1570
rect 3990 1550 4965 1565
rect 4990 1550 5000 1570
rect 5105 1570 5150 1580
rect 3000 1545 5000 1550
rect 5050 1500 5070 1560
rect 5105 1550 5115 1570
rect 5140 1565 5150 1570
rect 6385 1570 6430 1580
rect 6385 1565 6395 1570
rect 5140 1550 6395 1565
rect 6420 1565 6430 1570
rect 7230 1570 7275 1580
rect 7230 1565 7240 1570
rect 6420 1550 7240 1565
rect 7265 1565 7275 1570
rect 8510 1570 8555 1580
rect 8510 1565 8520 1570
rect 7265 1550 8520 1565
rect 8545 1550 8555 1570
rect 8660 1570 8705 1580
rect 5105 1545 8555 1550
rect 8590 1500 8610 1560
rect 8660 1550 8670 1570
rect 8695 1565 8705 1570
rect 9660 1570 9705 1580
rect 9660 1565 9670 1570
rect 8695 1550 9670 1565
rect 9695 1565 9705 1570
rect 10615 1570 10660 1580
rect 10615 1565 10625 1570
rect 9695 1550 10625 1565
rect 10650 1550 10660 1570
rect 10765 1570 10810 1580
rect 8660 1545 10660 1550
rect 10700 1500 10720 1560
rect 10765 1550 10775 1570
rect 10800 1565 10810 1570
rect 12090 1570 12135 1580
rect 12090 1565 12100 1570
rect 10800 1550 12100 1565
rect 12125 1550 12135 1570
rect 10765 1545 12135 1550
rect 33795 1545 33815 2315
rect 21725 1525 33815 1545
rect 12895 1500 12915 1510
rect -2425 1490 -835 1500
rect -2425 920 -2415 1490
rect -1645 920 -1615 1490
rect -845 920 -835 1490
rect -2425 910 -835 920
rect -25 1490 765 1500
rect -25 920 -15 1490
rect 755 920 765 1490
rect -25 910 765 920
rect 1575 1490 2365 1500
rect 1575 920 1585 1490
rect 2355 920 2365 1490
rect 1575 910 2365 920
rect 2405 1490 3195 1500
rect 2405 920 2415 1490
rect 3185 920 3195 1490
rect 2405 910 3195 920
rect 4005 1490 4795 1500
rect 4005 920 4015 1490
rect 4785 920 4795 1490
rect 4005 910 4795 920
rect 4835 1490 5625 1500
rect 4835 920 4845 1490
rect 5615 920 5625 1490
rect 4835 910 5625 920
rect 6435 1490 7225 1500
rect 6435 920 6445 1490
rect 7215 920 7225 1490
rect 6435 910 7225 920
rect 8035 1490 8825 1500
rect 8035 920 8045 1490
rect 8815 920 8825 1490
rect 8035 910 8825 920
rect 8865 1490 9655 1500
rect 8865 920 8875 1490
rect 9645 920 9655 1490
rect 8865 910 9655 920
rect 10465 1490 11255 1500
rect 10465 920 10475 1490
rect 11245 920 11255 1490
rect 10465 910 11255 920
rect 11295 1490 12085 1500
rect 11295 920 11305 1490
rect 12075 920 12085 1490
rect 11295 910 12085 920
rect 12895 1490 13685 1500
rect 12895 920 12905 1490
rect 13675 920 13685 1490
rect 21625 1485 21670 1495
rect 21625 1465 21635 1485
rect 21660 1465 21670 1485
rect 21625 1460 21670 1465
rect 21625 1445 21650 1460
rect 12895 910 13685 920
rect 16095 1425 21650 1445
rect 16095 1400 16115 1425
rect 18525 1400 18545 1425
rect 21725 1400 21745 1525
rect 21830 1485 21875 1495
rect 21830 1465 21840 1485
rect 21865 1465 21875 1485
rect 21830 1460 21875 1465
rect 21845 1445 21875 1460
rect 33840 1445 33860 2440
rect 33885 2400 33930 2410
rect 33885 2380 33895 2400
rect 33920 2395 33930 2400
rect 33920 2380 33945 2395
rect 33885 2375 33945 2380
rect 21845 1425 33860 1445
rect 25695 1400 25715 1425
rect 28125 1400 28145 1425
rect 16095 1390 16885 1400
rect 1635 840 1655 910
rect 4485 840 4505 910
rect 6745 845 6790 855
rect 6745 840 6755 845
rect 1635 825 6755 840
rect 6780 825 6790 845
rect 1635 820 6790 825
rect 6745 780 6790 790
rect 6745 775 6755 780
rect -3200 760 6755 775
rect 6780 760 6790 780
rect -3200 755 6790 760
rect 6460 720 6505 730
rect 6460 715 6470 720
rect 5665 700 6470 715
rect 6495 715 6505 720
rect 6745 720 6790 730
rect 6745 715 6755 720
rect 6495 700 6755 715
rect 6780 700 6790 720
rect 5665 695 6790 700
rect 0 665 45 675
rect 0 645 10 665
rect 35 660 45 665
rect 2430 665 2475 675
rect 2430 660 2440 665
rect 35 645 2440 660
rect 2465 660 2475 665
rect 4030 665 4075 675
rect 4030 660 4040 665
rect 2465 645 4040 660
rect 4065 660 4075 665
rect 5590 665 5635 675
rect 5590 660 5600 665
rect 4065 645 5600 660
rect 5625 645 5635 665
rect 0 640 5635 645
rect 4835 595 4855 640
rect 5665 595 5685 695
rect 5740 665 5785 675
rect 5740 645 5750 665
rect 5775 660 5785 665
rect 6840 660 6860 910
rect 6930 845 6975 855
rect 6930 825 6940 845
rect 6965 840 6975 845
rect 9155 840 9175 910
rect 12005 840 12025 910
rect 6965 825 12025 840
rect 6930 820 12025 825
rect 16095 820 16105 1390
rect 16875 820 16885 1390
rect 6930 780 6975 790
rect 6930 760 6940 780
rect 6965 775 6975 780
rect 9050 780 9095 790
rect 9050 775 9060 780
rect 6965 760 9060 775
rect 9085 760 9095 780
rect 6930 755 9095 760
rect 6930 720 6975 730
rect 6930 700 6940 720
rect 6965 715 6975 720
rect 9155 715 9175 820
rect 16095 810 16885 820
rect 17695 1390 18485 1400
rect 17695 820 17705 1390
rect 18475 820 18485 1390
rect 17695 810 18485 820
rect 18525 1390 19315 1400
rect 18525 820 18535 1390
rect 19305 820 19315 1390
rect 18525 810 19315 820
rect 20125 1390 20915 1400
rect 20125 820 20135 1390
rect 20905 820 20915 1390
rect 20125 810 20915 820
rect 21725 1390 22515 1400
rect 21725 820 21735 1390
rect 22505 820 22515 1390
rect 21725 810 22515 820
rect 23325 1390 24115 1400
rect 23325 820 23335 1390
rect 24105 820 24115 1390
rect 23325 810 24115 820
rect 24925 1390 25715 1400
rect 24925 820 24935 1390
rect 25705 820 25715 1390
rect 24925 810 25715 820
rect 25755 1390 26545 1400
rect 25755 820 25765 1390
rect 26535 820 26545 1390
rect 25755 810 26545 820
rect 27355 1390 28145 1400
rect 27355 820 27365 1390
rect 28135 820 28145 1390
rect 27355 810 28145 820
rect 28955 1390 30545 1400
rect 28955 820 28965 1390
rect 29735 820 29765 1390
rect 30535 820 30545 1390
rect 28955 810 30545 820
rect 28955 790 28975 810
rect 9215 780 9260 790
rect 9215 760 9225 780
rect 9250 775 9260 780
rect 16890 785 16935 790
rect 16890 775 16900 785
rect 9250 765 16900 775
rect 16925 775 16935 785
rect 19320 785 19365 790
rect 19320 775 19330 785
rect 16925 765 19330 775
rect 19355 775 19365 785
rect 20920 785 20965 790
rect 20920 775 20930 785
rect 19355 765 20930 775
rect 20955 775 20965 785
rect 23275 785 23320 790
rect 23275 775 23285 785
rect 20955 765 23285 775
rect 23310 775 23320 785
rect 24875 785 24920 790
rect 24875 775 24885 785
rect 23310 765 24885 775
rect 24910 775 24920 785
rect 27305 785 27350 790
rect 27305 775 27315 785
rect 24910 765 27315 775
rect 27340 765 27350 785
rect 9250 760 27350 765
rect 9215 755 27350 760
rect 28880 785 28975 790
rect 28880 765 28890 785
rect 28915 770 28975 785
rect 28915 765 28925 770
rect 28880 755 28925 765
rect 10490 720 10535 730
rect 10490 715 10500 720
rect 6965 700 10500 715
rect 10525 715 10535 720
rect 19245 720 19290 730
rect 19245 715 19255 720
rect 10525 700 19255 715
rect 19280 715 19290 720
rect 23275 720 23320 730
rect 23275 715 23285 720
rect 19280 700 23285 715
rect 23310 715 23320 720
rect 23310 700 33980 715
rect 6930 695 33980 700
rect 8060 665 8105 675
rect 8060 660 8070 665
rect 5775 645 8070 660
rect 8095 660 8105 665
rect 9620 665 9665 675
rect 9620 660 9630 665
rect 8095 645 9630 660
rect 9655 645 9665 665
rect 5740 640 9665 645
rect 8865 595 8885 640
rect 9695 595 9715 695
rect 9770 665 9815 675
rect 9770 645 9780 665
rect 9805 660 9815 665
rect 12090 665 12135 675
rect 12090 660 12100 665
rect 9805 645 12100 660
rect 12125 660 12135 665
rect 13690 665 13735 675
rect 13690 660 13700 665
rect 12125 645 13700 660
rect 13725 660 13735 665
rect 16045 665 16090 675
rect 16045 660 16055 665
rect 13725 645 16055 660
rect 16080 660 16090 665
rect 17645 665 17690 675
rect 17645 660 17655 665
rect 16080 645 17655 660
rect 17680 660 17690 665
rect 19965 665 20010 675
rect 19965 660 19975 665
rect 17680 645 19975 660
rect 20000 645 20010 665
rect 9770 640 20010 645
rect 12895 595 12915 640
rect 16865 595 16885 640
rect 20065 595 20085 695
rect 20115 665 20160 675
rect 20115 645 20125 665
rect 20150 660 20160 665
rect 21675 665 21720 675
rect 21675 660 21685 665
rect 20150 645 21685 660
rect 21710 660 21720 665
rect 23995 665 24040 675
rect 23995 660 24005 665
rect 21710 645 24005 660
rect 24030 645 24040 665
rect 20115 640 24040 645
rect 20895 595 20915 640
rect 24095 595 24115 695
rect 24145 665 24190 675
rect 24145 645 24155 665
rect 24180 660 24190 665
rect 25705 665 25750 675
rect 25705 660 25715 665
rect 24180 645 25715 660
rect 25740 660 25750 665
rect 27305 665 27350 675
rect 27305 660 27315 665
rect 25740 645 27315 660
rect 27340 660 27350 665
rect 29735 665 29780 675
rect 29735 660 29745 665
rect 27340 645 29745 660
rect 29770 645 29780 665
rect 24145 640 29780 645
rect 24925 595 24945 640
rect -3195 585 -1605 595
rect -3195 15 -3185 585
rect -2415 15 -2385 585
rect -1615 15 -1605 585
rect -3195 5 -1605 15
rect -795 585 -5 595
rect -795 15 -785 585
rect -15 15 -5 585
rect -795 5 -5 15
rect 805 585 1595 595
rect 805 15 815 585
rect 1585 15 1595 585
rect 805 5 1595 15
rect 1635 585 2425 595
rect 1635 15 1645 585
rect 2415 15 2425 585
rect 1635 5 2425 15
rect 3235 585 4025 595
rect 3235 15 3245 585
rect 4015 15 4025 585
rect 3235 5 4025 15
rect 4835 585 5625 595
rect 4835 15 4845 585
rect 5615 15 5625 585
rect 4835 5 5625 15
rect 5665 585 6455 595
rect 5665 15 5675 585
rect 6445 15 6455 585
rect 5665 5 6455 15
rect 7265 585 8055 595
rect 7265 15 7275 585
rect 8045 15 8055 585
rect 7265 5 8055 15
rect 8865 585 9655 595
rect 8865 15 8875 585
rect 9645 15 9655 585
rect 8865 5 9655 15
rect 9695 585 10485 595
rect 9695 15 9705 585
rect 10475 15 10485 585
rect 9695 5 10485 15
rect 11295 585 12085 595
rect 11295 15 11305 585
rect 12075 15 12085 585
rect 11295 5 12085 15
rect 12895 585 13685 595
rect 12895 15 12905 585
rect 13675 15 13685 585
rect 12895 5 13685 15
rect 14495 585 15285 595
rect 14495 15 14505 585
rect 15275 15 15285 585
rect 14495 5 15285 15
rect 16095 585 16885 595
rect 16095 15 16105 585
rect 16875 15 16885 585
rect 16095 5 16885 15
rect 17695 585 18485 595
rect 17695 15 17705 585
rect 18475 15 18485 585
rect 17695 5 18485 15
rect 19295 585 20085 595
rect 19295 15 19305 585
rect 20075 15 20085 585
rect 19295 5 20085 15
rect 20125 585 20915 595
rect 20125 15 20135 585
rect 20905 15 20915 585
rect 20125 5 20915 15
rect 21725 585 22515 595
rect 21725 15 21735 585
rect 22505 15 22515 585
rect 21725 5 22515 15
rect 23325 585 24115 595
rect 23325 15 23335 585
rect 24105 15 24115 585
rect 23325 5 24115 15
rect 24155 585 24945 595
rect 24155 15 24165 585
rect 24935 15 24945 585
rect 24155 5 24945 15
rect 25755 585 26545 595
rect 25755 15 25765 585
rect 26535 15 26545 585
rect 25755 5 26545 15
rect 27355 585 28145 595
rect 27355 15 27365 585
rect 28135 15 28145 585
rect 27355 5 28145 15
rect 28185 585 28975 595
rect 28185 15 28195 585
rect 28965 15 28975 585
rect 28185 5 28975 15
rect 29785 585 30575 595
rect 29785 15 29795 585
rect 30565 15 30575 585
rect 29785 5 30575 15
rect 31385 585 32975 595
rect 31385 15 31395 585
rect 32165 15 32195 585
rect 32965 15 32975 585
rect 31385 5 32975 15
rect -1625 -15 -1605 5
rect 805 -15 825 5
rect 3235 -15 3255 5
rect 7265 -15 7285 5
rect 11295 -15 11315 5
rect 14495 -15 14515 5
rect 18465 -15 18485 5
rect 22495 -15 22515 5
rect 26525 -15 26545 5
rect 28955 -15 28975 5
rect 31385 -15 31405 5
rect -1625 -20 -1555 -15
rect -1625 -35 -1590 -20
rect -1600 -40 -1590 -35
rect -1565 -40 -1555 -20
rect 805 -35 28975 -15
rect 31335 -20 31405 -15
rect -1600 -50 -1555 -40
rect 31335 -40 31345 -20
rect 31370 -35 31405 -20
rect 31370 -40 31380 -35
rect 31335 -50 31380 -40
<< viali >>
rect -2415 1690 -1645 2260
rect -1615 1690 -845 2260
rect -15 1690 755 2260
rect 2415 1690 3185 2260
rect 28135 1690 28905 2260
rect 30565 1690 31335 2260
rect 32165 1690 32935 2260
rect 32965 1690 33735 2260
rect -2415 920 -1645 1490
rect -1615 920 -845 1490
rect -15 920 755 1490
rect 2415 920 3185 1490
rect 4845 920 5615 1490
rect 8045 920 8815 1490
rect 10475 920 11245 1490
rect 12905 920 13675 1490
rect 17705 820 18475 1390
rect 20135 820 20905 1390
rect 23335 820 24105 1390
rect 25765 820 26535 1390
rect 28965 820 29735 1390
rect 29765 820 30535 1390
rect -3185 15 -2415 585
rect -2385 15 -1615 585
rect -785 15 -15 585
rect 1645 15 2415 585
rect 27365 15 28135 585
rect 29795 15 30565 585
rect 31395 15 32165 585
rect 32195 15 32965 585
<< metal1 >>
rect -2460 2260 33780 2275
rect -2460 1690 -2415 2260
rect -1645 1690 -1615 2260
rect -845 1690 -15 2260
rect 755 1690 2415 2260
rect 3185 1690 28135 2260
rect 28905 1690 30565 2260
rect 31335 1690 32165 2260
rect 32935 1690 32965 2260
rect 33735 1690 33780 2260
rect -2460 1675 33780 1690
rect -2460 1490 13725 1675
rect 17595 1640 33780 1675
rect -2460 920 -2415 1490
rect -1645 920 -1615 1490
rect -845 920 -15 1490
rect 755 920 2415 1490
rect 3185 920 4845 1490
rect 5615 920 8045 1490
rect 8815 920 10475 1490
rect 11245 920 12905 1490
rect 13675 920 13725 1490
rect -2460 905 13725 920
rect 16090 1390 30550 1405
rect 16090 820 17705 1390
rect 18475 820 20135 1390
rect 20905 820 23335 1390
rect 24105 820 25765 1390
rect 26535 820 28965 1390
rect 29735 820 29765 1390
rect 30535 820 30550 1390
rect 16090 600 30550 820
rect -3200 585 32980 600
rect -3200 15 -3185 585
rect -2415 15 -2385 585
rect -1615 15 -785 585
rect -15 15 1645 585
rect 2415 15 27365 585
rect 28135 15 29795 585
rect 30565 15 31395 585
rect 32165 15 32195 585
rect 32965 15 32980 585
rect -3200 0 32980 15
<< labels >>
rlabel locali -3230 1615 -3230 1615 7 Vbp
port 1 w
rlabel locali -3200 765 -3200 765 7 Vbn
port 2 w
rlabel locali 33945 2450 33945 2450 3 Vcp
port 3 e
rlabel locali 33980 705 33980 705 3 Vcn
port 4 e
rlabel metal1 -3200 595 -3200 595 7 VN
port 5 w
rlabel metal1 -2460 910 -2460 910 7 VP
port 6 w
<< end >>
