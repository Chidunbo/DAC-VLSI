magic
tech sky130A
timestamp 1693780072
<< nwell >>
rect -240 45 -30 185
<< nmos >>
rect -120 -90 -105 10
<< pmos >>
rect -120 65 -105 165
<< ndiff >>
rect -170 -5 -120 10
rect -170 -75 -155 -5
rect -135 -75 -120 -5
rect -170 -90 -120 -75
rect -105 -5 -55 10
rect -105 -75 -90 -5
rect -70 -75 -55 -5
rect -105 -90 -55 -75
<< pdiff >>
rect -170 150 -120 165
rect -170 80 -155 150
rect -135 80 -120 150
rect -170 65 -120 80
rect -105 150 -55 165
rect -105 80 -90 150
rect -70 80 -55 150
rect -105 65 -55 80
<< ndiffc >>
rect -155 -75 -135 -5
rect -90 -75 -70 -5
<< pdiffc >>
rect -155 80 -135 150
rect -90 80 -70 150
<< psubdiff >>
rect -220 -5 -170 10
rect -220 -75 -205 -5
rect -185 -75 -170 -5
rect -220 -90 -170 -75
<< nsubdiff >>
rect -220 150 -170 165
rect -220 80 -205 150
rect -185 80 -170 150
rect -220 65 -170 80
<< psubdiffcont >>
rect -205 -75 -185 -5
<< nsubdiffcont >>
rect -205 80 -185 150
<< poly >>
rect -120 165 -105 180
rect -120 10 -105 65
rect -120 -105 -105 -90
rect -145 -115 -105 -105
rect -145 -135 -135 -115
rect -115 -135 -105 -115
rect -145 -145 -105 -135
<< polycont >>
rect -135 -135 -115 -115
<< locali >>
rect -215 150 -125 160
rect -215 80 -205 150
rect -185 80 -155 150
rect -135 80 -125 150
rect -215 70 -125 80
rect -100 150 -60 160
rect -100 80 -90 150
rect -70 80 -60 150
rect -100 70 -60 80
rect -80 5 -60 70
rect -215 -5 -125 5
rect -215 -75 -205 -5
rect -185 -75 -155 -5
rect -135 -75 -125 -5
rect -215 -85 -125 -75
rect -100 -5 -60 5
rect -100 -75 -90 -5
rect -70 -75 -60 -5
rect -100 -85 -60 -75
rect -80 -105 -60 -85
rect -240 -115 -105 -105
rect -240 -125 -135 -115
rect -145 -135 -135 -125
rect -115 -135 -105 -115
rect -80 -125 -30 -105
rect -145 -145 -105 -135
<< viali >>
rect -205 80 -185 150
rect -155 80 -135 150
rect -205 -75 -185 -5
rect -155 -75 -135 -5
<< metal1 >>
rect -240 150 -30 160
rect -240 80 -205 150
rect -185 80 -155 150
rect -135 80 -30 150
rect -240 70 -30 80
rect -240 -5 -30 5
rect -240 -75 -205 -5
rect -185 -75 -155 -5
rect -135 -75 -30 -5
rect -240 -85 -30 -75
<< labels >>
rlabel locali -240 -115 -240 -115 7 A
port 1 w
rlabel locali -30 -115 -30 -115 3 Y
port 2 e
rlabel metal1 -240 115 -240 115 7 VP
port 3 w
rlabel metal1 -240 -40 -240 -40 7 VN
port 4 w
<< end >>
