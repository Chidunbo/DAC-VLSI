magic
tech sky130A
timestamp 1700362378
<< nwell >>
rect -1790 4695 18445 8265
<< nmos >>
rect -930 3350 -130 4550
rect 670 3350 1470 4550
rect 3100 3350 3900 4550
rect 4700 3350 5500 4550
rect 7125 3350 7925 4550
rect 8725 3350 9525 4550
rect 11150 3350 11950 4550
rect 12750 3350 13550 4550
rect 15180 3350 15980 4550
rect 16780 3350 17580 4550
rect 725 1155 1525 2355
rect 2325 1155 3125 2355
rect 3925 1155 4725 2355
rect 5525 1155 6325 2355
rect 7125 1155 7925 2355
rect 8725 1155 9525 2355
rect 10325 1155 11125 2355
rect 11925 1155 12725 2355
rect 13525 1155 14325 2355
rect 15125 1155 15925 2355
<< pmos >>
rect 725 6950 1525 8150
rect 2325 6950 3125 8150
rect 3925 6950 4725 8150
rect 5525 6950 6325 8150
rect 7125 6950 7925 8150
rect 8725 6950 9525 8150
rect 10325 6950 11125 8150
rect 11925 6950 12725 8150
rect 13525 6950 14325 8150
rect 15125 6950 15925 8150
rect -930 4755 -130 5955
rect 670 4755 1470 5955
rect 3100 4755 3900 5955
rect 4700 4755 5500 5955
rect 7125 4755 7925 5955
rect 8725 4755 9525 5955
rect 11150 4755 11950 5955
rect 12750 4755 13550 5955
rect 15180 4755 15980 5955
rect 16780 4755 17580 5955
<< ndiff >>
rect -1730 4535 -930 4550
rect -1730 3365 -1715 4535
rect -945 3365 -930 4535
rect -1730 3350 -930 3365
rect -130 4535 670 4550
rect -130 3365 -115 4535
rect 655 3365 670 4535
rect -130 3350 670 3365
rect 1470 4535 2270 4550
rect 1470 3365 1485 4535
rect 2255 3365 2270 4535
rect 1470 3350 2270 3365
rect 2300 4535 3100 4550
rect 2300 3365 2315 4535
rect 3085 3365 3100 4535
rect 2300 3350 3100 3365
rect 3900 4535 4700 4550
rect 3900 3365 3915 4535
rect 4685 3365 4700 4535
rect 3900 3350 4700 3365
rect 5500 4535 6300 4550
rect 5500 3365 5515 4535
rect 6285 3365 6300 4535
rect 5500 3350 6300 3365
rect 6330 4535 7125 4550
rect 6330 3365 6345 4535
rect 7115 3365 7125 4535
rect 6330 3350 7125 3365
rect 7925 4535 8725 4550
rect 7925 3365 7940 4535
rect 8710 3365 8725 4535
rect 7925 3350 8725 3365
rect 9525 4535 10320 4550
rect 9525 3365 9535 4535
rect 10305 3365 10320 4535
rect 9525 3350 10320 3365
rect 10350 4535 11150 4550
rect 10350 3365 10365 4535
rect 11135 3365 11150 4535
rect 10350 3350 11150 3365
rect 11950 4535 12750 4550
rect 11950 3365 11965 4535
rect 12735 3365 12750 4535
rect 11950 3350 12750 3365
rect 13550 4535 14350 4550
rect 13550 3365 13565 4535
rect 14335 3365 14350 4535
rect 13550 3350 14350 3365
rect 14380 4535 15180 4550
rect 14380 3365 14395 4535
rect 15165 3365 15180 4535
rect 14380 3350 15180 3365
rect 15980 4535 16780 4550
rect 15980 3365 15995 4535
rect 16765 3365 16780 4535
rect 15980 3350 16780 3365
rect 17580 4535 18380 4550
rect 17580 3365 17595 4535
rect 18365 3365 18380 4535
rect 17580 3350 18380 3365
rect -75 2340 725 2355
rect -75 1170 -60 2340
rect 710 1170 725 2340
rect -75 1155 725 1170
rect 1525 2340 2325 2355
rect 1525 1170 1540 2340
rect 2310 1170 2325 2340
rect 1525 1155 2325 1170
rect 3125 2340 3925 2355
rect 3125 1170 3140 2340
rect 3910 1170 3925 2340
rect 3125 1155 3925 1170
rect 4725 2340 5525 2355
rect 4725 1170 4740 2340
rect 5510 1170 5525 2340
rect 4725 1155 5525 1170
rect 6325 2340 7125 2355
rect 6325 1170 6340 2340
rect 7110 1170 7125 2340
rect 6325 1155 7125 1170
rect 7925 2340 8725 2355
rect 7925 1170 7940 2340
rect 8710 1170 8725 2340
rect 7925 1155 8725 1170
rect 9525 2340 10325 2355
rect 9525 1170 9540 2340
rect 10310 1170 10325 2340
rect 9525 1155 10325 1170
rect 11125 2340 11925 2355
rect 11125 1170 11140 2340
rect 11910 1170 11925 2340
rect 11125 1155 11925 1170
rect 12725 2340 13525 2355
rect 12725 1170 12740 2340
rect 13510 1170 13525 2340
rect 12725 1155 13525 1170
rect 14325 2340 15125 2355
rect 14325 1170 14340 2340
rect 15110 1170 15125 2340
rect 14325 1155 15125 1170
rect 15925 2340 16725 2355
rect 15925 1170 15940 2340
rect 16710 1170 16725 2340
rect 15925 1155 16725 1170
<< pdiff >>
rect -75 8135 725 8150
rect -75 6965 -60 8135
rect 710 6965 725 8135
rect -75 6950 725 6965
rect 1525 8135 2325 8150
rect 1525 6965 1540 8135
rect 2310 6965 2325 8135
rect 1525 6950 2325 6965
rect 3125 8135 3925 8150
rect 3125 6965 3140 8135
rect 3910 6965 3925 8135
rect 3125 6950 3925 6965
rect 4725 8135 5525 8150
rect 4725 6965 4740 8135
rect 5510 6965 5525 8135
rect 4725 6950 5525 6965
rect 6325 8135 7125 8150
rect 6325 6965 6340 8135
rect 7110 6965 7125 8135
rect 6325 6950 7125 6965
rect 7925 8135 8725 8150
rect 7925 6965 7940 8135
rect 8710 6965 8725 8135
rect 7925 6950 8725 6965
rect 9525 8135 10325 8150
rect 9525 6965 9540 8135
rect 10310 6965 10325 8135
rect 9525 6950 10325 6965
rect 11125 8135 11925 8150
rect 11125 6965 11140 8135
rect 11910 6965 11925 8135
rect 11125 6950 11925 6965
rect 12725 8135 13525 8150
rect 12725 6965 12740 8135
rect 13510 6965 13525 8135
rect 12725 6950 13525 6965
rect 14325 8135 15125 8150
rect 14325 6965 14340 8135
rect 15110 6965 15125 8135
rect 14325 6950 15125 6965
rect 15925 8135 16725 8150
rect 15925 6965 15940 8135
rect 16710 6965 16725 8135
rect 15925 6950 16725 6965
rect -1730 5940 -930 5955
rect -1730 4770 -1715 5940
rect -945 4770 -930 5940
rect -1730 4755 -930 4770
rect -130 5940 670 5955
rect -130 4770 -115 5940
rect 655 4770 670 5940
rect -130 4755 670 4770
rect 1470 5940 2270 5955
rect 1470 4770 1485 5940
rect 2255 4770 2270 5940
rect 1470 4755 2270 4770
rect 2300 5940 3100 5955
rect 2300 4770 2315 5940
rect 3085 4770 3100 5940
rect 2300 4755 3100 4770
rect 3900 5940 4700 5955
rect 3900 4770 3915 5940
rect 4685 4770 4700 5940
rect 3900 4755 4700 4770
rect 5500 5940 6300 5955
rect 5500 4770 5515 5940
rect 6285 4770 6300 5940
rect 5500 4755 6300 4770
rect 6330 5940 7125 5955
rect 6330 4770 6345 5940
rect 7115 4770 7125 5940
rect 6330 4755 7125 4770
rect 7925 5940 8725 5955
rect 7925 4770 7940 5940
rect 8710 4770 8725 5940
rect 7925 4755 8725 4770
rect 9525 5940 10320 5955
rect 9525 4770 9535 5940
rect 10305 4770 10320 5940
rect 9525 4755 10320 4770
rect 10350 5940 11150 5955
rect 10350 4770 10365 5940
rect 11135 4770 11150 5940
rect 10350 4755 11150 4770
rect 11950 5940 12750 5955
rect 11950 4770 11965 5940
rect 12735 4770 12750 5940
rect 11950 4755 12750 4770
rect 13550 5940 14350 5955
rect 13550 4770 13565 5940
rect 14335 4770 14350 5940
rect 13550 4755 14350 4770
rect 14380 5940 15180 5955
rect 14380 4770 14395 5940
rect 15165 4770 15180 5940
rect 14380 4755 15180 4770
rect 15980 5940 16780 5955
rect 15980 4770 15995 5940
rect 16765 4770 16780 5940
rect 15980 4755 16780 4770
rect 17580 5940 18380 5955
rect 17580 4770 17595 5940
rect 18365 4770 18380 5940
rect 17580 4755 18380 4770
<< ndiffc >>
rect -1715 3365 -945 4535
rect -115 3365 655 4535
rect 1485 3365 2255 4535
rect 2315 3365 3085 4535
rect 3915 3365 4685 4535
rect 5515 3365 6285 4535
rect 6345 3365 7115 4535
rect 7940 3365 8710 4535
rect 9535 3365 10305 4535
rect 10365 3365 11135 4535
rect 11965 3365 12735 4535
rect 13565 3365 14335 4535
rect 14395 3365 15165 4535
rect 15995 3365 16765 4535
rect 17595 3365 18365 4535
rect -60 1170 710 2340
rect 1540 1170 2310 2340
rect 3140 1170 3910 2340
rect 4740 1170 5510 2340
rect 6340 1170 7110 2340
rect 7940 1170 8710 2340
rect 9540 1170 10310 2340
rect 11140 1170 11910 2340
rect 12740 1170 13510 2340
rect 14340 1170 15110 2340
rect 15940 1170 16710 2340
<< pdiffc >>
rect -60 6965 710 8135
rect 1540 6965 2310 8135
rect 3140 6965 3910 8135
rect 4740 6965 5510 8135
rect 6340 6965 7110 8135
rect 7940 6965 8710 8135
rect 9540 6965 10310 8135
rect 11140 6965 11910 8135
rect 12740 6965 13510 8135
rect 14340 6965 15110 8135
rect 15940 6965 16710 8135
rect -1715 4770 -945 5940
rect -115 4770 655 5940
rect 1485 4770 2255 5940
rect 2315 4770 3085 5940
rect 3915 4770 4685 5940
rect 5515 4770 6285 5940
rect 6345 4770 7115 5940
rect 7940 4770 8710 5940
rect 9535 4770 10305 5940
rect 10365 4770 11135 5940
rect 11965 4770 12735 5940
rect 13565 4770 14335 5940
rect 14395 4770 15165 5940
rect 15995 4770 16765 5940
rect 17595 4770 18365 5940
<< psubdiff >>
rect 2340 3250 3540 3265
rect -825 3225 375 3240
rect -825 2505 -810 3225
rect 360 2505 375 3225
rect -825 2490 375 2505
rect 2340 2530 2355 3250
rect 3525 2530 3540 3250
rect 2340 2515 3540 2530
rect 6385 3240 7585 3255
rect 6385 2520 6400 3240
rect 7570 2520 7585 3240
rect 6385 2505 7585 2520
rect 9065 3240 10265 3255
rect 9065 2520 9080 3240
rect 10250 2520 10265 3240
rect 13110 3250 14310 3265
rect 13110 2530 13125 3250
rect 14295 2530 14310 3250
rect 9065 2505 10265 2520
rect 13110 2515 14310 2530
rect 16275 3225 17475 3240
rect 16275 2505 16290 3225
rect 17460 2505 17475 3225
rect 16275 2490 17475 2505
<< nsubdiff >>
rect -825 6800 375 6815
rect -825 6080 -810 6800
rect 360 6080 375 6800
rect -825 6065 375 6080
rect 2340 6775 3540 6790
rect 6385 6785 7585 6800
rect 2340 6055 2355 6775
rect 3525 6055 3540 6775
rect 2340 6040 3540 6055
rect 6385 6065 6400 6785
rect 7570 6065 7585 6785
rect 6385 6050 7585 6065
rect 9065 6785 10265 6800
rect 16275 6800 17475 6815
rect 9065 6065 9080 6785
rect 10250 6065 10265 6785
rect 9065 6050 10265 6065
rect 13110 6775 14310 6790
rect 13110 6055 13125 6775
rect 14295 6055 14310 6775
rect 16275 6080 16290 6800
rect 17460 6080 17475 6800
rect 16275 6065 17475 6080
rect 13110 6040 14310 6055
<< psubdiffcont >>
rect -810 2505 360 3225
rect 2355 2530 3525 3250
rect 6400 2520 7570 3240
rect 9080 2520 10250 3240
rect 13125 2530 14295 3250
rect 16290 2505 17460 3225
<< nsubdiffcont >>
rect -810 6080 360 6800
rect 2355 6055 3525 6775
rect 6400 6065 7570 6785
rect 9080 6065 10250 6785
rect 13125 6055 14295 6775
rect 16290 6080 17460 6800
<< poly >>
rect 725 8205 1525 8215
rect 725 8185 735 8205
rect 1515 8185 1525 8205
rect 725 8150 1525 8185
rect 2325 8200 14325 8225
rect 2325 8150 3125 8200
rect 3925 8150 4725 8200
rect 5525 8150 6325 8175
rect 7125 8150 7925 8200
rect 8725 8150 9525 8200
rect 10325 8150 11125 8175
rect 11925 8150 12725 8200
rect 13525 8150 14325 8200
rect 15125 8205 15925 8215
rect 15125 8185 15135 8205
rect 15915 8185 15925 8205
rect 15125 8150 15925 8185
rect 725 6925 1525 6950
rect 2325 6895 3125 6950
rect 3925 6920 4725 6950
rect -1790 6870 3125 6895
rect 5525 6915 6325 6950
rect 7125 6925 7925 6950
rect 8725 6925 9525 6950
rect 5525 6895 5535 6915
rect 6315 6895 6325 6915
rect 5525 6885 6325 6895
rect 10325 6915 11125 6950
rect 11925 6925 12725 6950
rect 13525 6925 14325 6950
rect 15125 6925 15925 6950
rect 10325 6895 10335 6915
rect 11115 6895 11125 6915
rect 10325 6885 11125 6895
rect 4790 6840 11860 6855
rect 4790 6800 4805 6840
rect 4845 6825 11805 6840
rect 4845 6800 4860 6825
rect 11790 6800 11805 6825
rect 11845 6800 11860 6840
rect 4790 6785 4860 6800
rect 11790 6785 11860 6800
rect -1790 6025 670 6035
rect -1790 6005 15980 6025
rect -930 5955 -130 5980
rect 670 5955 1470 6005
rect 3100 5955 3900 6005
rect 7125 6000 9525 6005
rect 4700 5955 5500 5980
rect 7125 5955 7925 6000
rect 8725 5955 9525 6000
rect 11150 5955 11950 5980
rect 12750 5955 13550 6005
rect 15180 5955 15980 6005
rect 16780 5955 17580 5980
rect -930 4720 -130 4755
rect 670 4730 1470 4755
rect 3100 4730 3900 4755
rect -930 4700 -920 4720
rect -140 4700 -130 4720
rect -930 4690 -130 4700
rect 4700 4720 5500 4755
rect 7125 4730 7925 4755
rect 8725 4730 9525 4755
rect 4700 4700 4710 4720
rect 5490 4700 5500 4720
rect 4700 4690 5500 4700
rect 11150 4720 11950 4755
rect 12750 4730 13550 4755
rect 15180 4730 15980 4755
rect 11150 4700 11160 4720
rect 11940 4700 11950 4720
rect 11150 4690 11950 4700
rect 16780 4720 17580 4755
rect 16780 4700 16790 4720
rect 17570 4700 17580 4720
rect 16780 4690 17580 4700
rect 9530 4650 18445 4665
rect 9530 4615 9545 4650
rect 10300 4640 18445 4650
rect 10300 4615 10315 4640
rect -930 4605 -130 4615
rect -930 4585 -920 4605
rect -140 4585 -130 4605
rect -930 4550 -130 4585
rect 4700 4605 5500 4615
rect 4700 4585 4710 4605
rect 5490 4585 5500 4605
rect 9530 4600 10315 4615
rect 11150 4605 11950 4615
rect 670 4550 1470 4575
rect 3100 4550 3900 4575
rect 4700 4550 5500 4585
rect 11150 4585 11160 4605
rect 11940 4585 11950 4605
rect 7125 4550 7925 4575
rect 8725 4550 9525 4575
rect 11150 4550 11950 4585
rect 16780 4605 17580 4615
rect 16780 4585 16790 4605
rect 17570 4585 17580 4605
rect 12750 4550 13550 4575
rect 15180 4550 15980 4575
rect 16780 4550 17580 4585
rect -930 3325 -130 3350
rect 670 3300 1470 3350
rect 3100 3300 3900 3350
rect 4700 3325 5500 3350
rect 7125 3305 7925 3350
rect 8725 3305 9525 3350
rect 11150 3325 11950 3350
rect 7125 3300 9525 3305
rect 12750 3300 13550 3350
rect 15180 3300 15980 3350
rect 16780 3325 17580 3350
rect -940 3280 15980 3300
rect -940 3270 670 3280
rect -940 3165 -910 3270
rect -1790 3135 -910 3165
rect 1510 3220 2325 3230
rect 1510 3200 1525 3220
rect 2305 3200 2325 3220
rect 1510 3190 2325 3200
rect -1790 2435 2210 2450
rect -1790 2420 2155 2435
rect 2140 2395 2155 2420
rect 2195 2395 2210 2435
rect 2140 2380 2210 2395
rect 2295 2420 2325 3190
rect 4790 2510 4860 2525
rect 4790 2475 4805 2510
rect 3390 2470 4805 2475
rect 4845 2480 4860 2510
rect 11790 2510 11860 2525
rect 14325 3220 15140 3230
rect 14325 3200 14345 3220
rect 15125 3200 15140 3220
rect 14325 3190 15140 3200
rect 11790 2480 11805 2510
rect 4845 2470 11805 2480
rect 11845 2470 11860 2510
rect 3390 2455 11860 2470
rect 3390 2450 4790 2455
rect 3390 2435 3460 2450
rect 2295 2380 3125 2420
rect 3390 2395 3405 2435
rect 3445 2395 3460 2435
rect 14325 2420 14355 3190
rect 3390 2380 3460 2395
rect 3925 2410 4725 2420
rect 3925 2390 3935 2410
rect 4715 2390 4725 2410
rect 725 2355 1525 2380
rect 2325 2355 3125 2380
rect 3925 2355 4725 2390
rect 5525 2410 6325 2420
rect 5525 2390 5535 2410
rect 6315 2390 6325 2410
rect 5525 2355 6325 2390
rect 10325 2410 11125 2420
rect 10325 2390 10335 2410
rect 11115 2390 11125 2410
rect 7125 2355 7925 2380
rect 8725 2355 9525 2380
rect 10325 2355 11125 2390
rect 11925 2410 12725 2420
rect 11925 2390 11935 2410
rect 12715 2390 12725 2410
rect 11925 2355 12725 2390
rect 13525 2380 14355 2420
rect 13525 2355 14325 2380
rect 15125 2355 15925 2380
rect 725 1120 1525 1155
rect 725 1100 735 1120
rect 1515 1100 1525 1120
rect 725 1090 1525 1100
rect 2325 1055 3125 1155
rect 3925 1105 4725 1155
rect 5525 1130 6325 1155
rect 7125 1105 7925 1155
rect 8725 1105 9525 1155
rect 10325 1130 11125 1155
rect 11925 1105 12725 1155
rect 3925 1080 12725 1105
rect 13525 1055 14325 1155
rect 15125 1120 15925 1155
rect 15125 1100 15135 1120
rect 15915 1100 15925 1120
rect 15125 1090 15925 1100
rect 2325 1030 14325 1055
<< polycont >>
rect 735 8185 1515 8205
rect 15135 8185 15915 8205
rect 5535 6895 6315 6915
rect 10335 6895 11115 6915
rect 4805 6800 4845 6840
rect 11805 6800 11845 6840
rect -920 4700 -140 4720
rect 4710 4700 5490 4720
rect 11160 4700 11940 4720
rect 16790 4700 17570 4720
rect 9545 4615 10300 4650
rect -920 4585 -140 4605
rect 4710 4585 5490 4605
rect 11160 4585 11940 4605
rect 16790 4585 17570 4605
rect 1525 3200 2305 3220
rect 2155 2395 2195 2435
rect 4805 2470 4845 2510
rect 14345 3200 15125 3220
rect 11805 2470 11845 2510
rect 3405 2395 3445 2435
rect 3935 2390 4715 2410
rect 5535 2390 6315 2410
rect 10335 2390 11115 2410
rect 11935 2390 12715 2410
rect 735 1100 1515 1120
rect 15135 1100 15915 1120
<< locali >>
rect 1690 8230 12415 8235
rect 725 8205 1525 8215
rect 725 8185 735 8205
rect 1515 8185 1525 8205
rect 725 8175 1525 8185
rect 1690 8190 14905 8230
rect 1690 8145 2320 8190
rect 14330 8145 14905 8190
rect 15125 8205 15925 8215
rect 15125 8185 15135 8205
rect 15915 8185 15925 8205
rect 15125 8175 15925 8185
rect -70 8135 720 8145
rect -70 6965 -60 8135
rect 710 6965 720 8135
rect -70 6955 720 6965
rect 1530 8135 2320 8145
rect 1530 6965 1540 8135
rect 2310 6965 2320 8135
rect 1530 6955 2320 6965
rect 3130 8135 3920 8145
rect 3130 6965 3140 8135
rect 3910 6965 3920 8135
rect 3130 6955 3920 6965
rect 4730 8135 5520 8145
rect 4730 6965 4740 8135
rect 5510 6965 5520 8135
rect 4730 6955 5520 6965
rect 6330 8135 7120 8145
rect 6330 6965 6340 8135
rect 7110 6965 7120 8135
rect 6330 6955 7120 6965
rect 7930 8135 8720 8145
rect 7930 6965 7940 8135
rect 8710 6965 8720 8135
rect 1530 6905 1790 6955
rect 550 6845 1790 6905
rect 4790 6905 5465 6955
rect 5525 6915 6325 6925
rect -820 6800 370 6810
rect -820 6080 -810 6800
rect 360 6080 370 6800
rect -820 6070 370 6080
rect 550 6045 620 6845
rect 4790 6840 4860 6905
rect 5525 6895 5535 6915
rect 6315 6895 6325 6915
rect 5525 6885 6325 6895
rect 4790 6800 4805 6840
rect 4845 6800 4860 6840
rect 2345 6775 3535 6785
rect 2345 6055 2355 6775
rect 3525 6055 3535 6775
rect 2345 6045 3535 6055
rect 4790 6050 4860 6800
rect 6390 6785 7580 6795
rect 6390 6065 6400 6785
rect 7570 6065 7580 6785
rect 6390 6055 7580 6065
rect -130 5950 620 6045
rect 3905 5985 4860 6050
rect -1725 5940 -935 5950
rect -1725 4770 -1715 5940
rect -945 4770 -935 5940
rect -1725 4760 -935 4770
rect -125 5940 665 5950
rect -125 4770 -115 5940
rect 655 4770 665 5940
rect -125 4760 665 4770
rect 1475 5940 2265 5950
rect 1475 4770 1485 5940
rect 2255 4770 2265 5940
rect -930 4720 -130 4730
rect -930 4700 -920 4720
rect -140 4700 -130 4720
rect -930 4690 -130 4700
rect -930 4605 -130 4615
rect -930 4585 -920 4605
rect -140 4585 -130 4605
rect -930 4575 -130 4585
rect -1725 4535 -935 4545
rect -1725 3365 -1715 4535
rect -945 3365 -935 4535
rect -1725 3355 -935 3365
rect -125 4535 665 4545
rect -125 3365 -115 4535
rect 655 3365 665 4535
rect -125 3355 665 3365
rect 1475 4535 2265 4770
rect 1475 3365 1485 4535
rect 2255 3365 2265 4535
rect 1475 3355 2265 3365
rect -130 3315 620 3355
rect -1790 3260 620 3315
rect -820 3225 370 3235
rect -820 2505 -810 3225
rect 360 2505 370 3225
rect -820 2495 370 2505
rect 550 2460 620 3260
rect 1510 3230 2265 3355
rect 2305 5940 3095 5950
rect 2305 4770 2315 5940
rect 3085 4770 3095 5940
rect 2305 4535 3095 4770
rect 3905 5940 4695 5985
rect 3905 4770 3915 5940
rect 4685 4770 4695 5940
rect 3905 4760 4695 4770
rect 5505 5940 6295 5950
rect 5505 4770 5515 5940
rect 6285 4770 6295 5940
rect 5505 4760 6295 4770
rect 6335 5940 7125 5950
rect 6335 4770 6345 5940
rect 7115 4770 7125 5940
rect 6335 4760 7125 4770
rect 7930 5940 8720 6965
rect 9530 8135 10320 8145
rect 9530 6965 9540 8135
rect 10310 6965 10320 8135
rect 9530 6955 10320 6965
rect 11130 8135 11920 8145
rect 11130 6965 11140 8135
rect 11910 6965 11920 8135
rect 11130 6955 11920 6965
rect 12730 8135 13520 8145
rect 12730 6965 12740 8135
rect 13510 6965 13520 8135
rect 12730 6955 13520 6965
rect 14330 8135 15120 8145
rect 14330 6965 14340 8135
rect 15110 6965 15120 8135
rect 10325 6915 11125 6925
rect 10325 6895 10335 6915
rect 11115 6895 11125 6915
rect 11185 6905 11860 6955
rect 10325 6885 11125 6895
rect 11790 6840 11860 6905
rect 14330 6905 15120 6965
rect 15930 8135 16720 8145
rect 15930 6965 15940 8135
rect 16710 6965 16720 8135
rect 15930 6955 16720 6965
rect 14330 6845 16055 6905
rect 11790 6800 11805 6840
rect 11845 6800 11860 6840
rect 9070 6785 10260 6795
rect 9070 6065 9080 6785
rect 10250 6065 10260 6785
rect 9070 6055 10260 6065
rect 11790 6050 11860 6800
rect 13115 6775 14305 6785
rect 13115 6055 13125 6775
rect 14295 6055 14305 6775
rect 11790 5985 12745 6050
rect 13115 6045 14305 6055
rect 7930 4770 7940 5940
rect 8710 4770 8720 5940
rect 7930 4760 8720 4770
rect 9525 5940 10315 5950
rect 9525 4770 9535 5940
rect 10305 4770 10315 5940
rect 9525 4760 10315 4770
rect 10355 5940 11145 5950
rect 10355 4770 10365 5940
rect 11135 4770 11145 5940
rect 10355 4760 11145 4770
rect 11955 5940 12745 5985
rect 15985 5990 16055 6845
rect 16280 6800 17470 6810
rect 16280 6080 16290 6800
rect 17460 6080 17470 6800
rect 16280 6070 17470 6080
rect 15985 5950 16780 5990
rect 11955 4770 11965 5940
rect 12735 4770 12745 5940
rect 11955 4760 12745 4770
rect 13555 5940 14345 5950
rect 13555 4770 13565 5940
rect 14335 4770 14345 5940
rect 4700 4720 5500 4730
rect 4700 4700 4710 4720
rect 5490 4700 5500 4720
rect 4700 4690 5500 4700
rect 6335 4685 7120 4760
rect 9530 4685 10315 4760
rect 11150 4720 11950 4730
rect 11150 4700 11160 4720
rect 11940 4700 11950 4720
rect 11150 4690 11950 4700
rect 6335 4650 10315 4685
rect 6335 4625 9545 4650
rect 4700 4605 5500 4615
rect 4700 4585 4710 4605
rect 5490 4585 5500 4605
rect 4700 4575 5500 4585
rect 6335 4545 7120 4625
rect 9530 4615 9545 4625
rect 10300 4615 10315 4650
rect 9530 4545 10315 4615
rect 11150 4605 11950 4615
rect 11150 4585 11160 4605
rect 11940 4585 11950 4605
rect 11150 4575 11950 4585
rect 2305 3365 2315 4535
rect 3085 3365 3095 4535
rect 2305 3355 3095 3365
rect 3905 4535 4695 4545
rect 3905 3365 3915 4535
rect 4685 3365 4695 4535
rect 2305 3315 3060 3355
rect 3905 3320 4695 3365
rect 5505 4535 6295 4545
rect 5505 3365 5515 4535
rect 6285 3365 6295 4535
rect 5505 3355 6295 3365
rect 6335 4535 7125 4545
rect 6335 3365 6345 4535
rect 7115 3365 7125 4535
rect 6335 3355 7125 3365
rect 7930 4535 8720 4545
rect 7930 3365 7940 4535
rect 8710 3365 8720 4535
rect 2305 3280 3615 3315
rect 2345 3250 3535 3260
rect 1510 3220 2325 3230
rect 1510 3200 1525 3220
rect 2305 3200 2325 3220
rect 1510 3190 2325 3200
rect 2345 2530 2355 3250
rect 3525 2530 3535 3250
rect 2345 2520 3535 2530
rect 550 2400 1790 2460
rect 1530 2350 1790 2400
rect 2140 2435 3460 2450
rect 2140 2395 2155 2435
rect 2195 2415 3405 2435
rect 2195 2395 2210 2415
rect 2140 2380 2210 2395
rect 3390 2395 3405 2415
rect 3445 2395 3460 2435
rect 3390 2380 3460 2395
rect 3575 2420 3615 3280
rect 3905 3255 4860 3320
rect 4790 2510 4860 3255
rect 6390 3240 7580 3250
rect 6390 2520 6400 3240
rect 7570 2520 7580 3240
rect 6390 2510 7580 2520
rect 4790 2470 4805 2510
rect 4845 2470 4860 2510
rect 3575 2410 4725 2420
rect 3575 2390 3935 2410
rect 4715 2390 4725 2410
rect 3575 2380 4725 2390
rect 4790 2400 4860 2470
rect 5525 2410 6325 2420
rect 4790 2350 5465 2400
rect 5525 2390 5535 2410
rect 6315 2390 6325 2410
rect 5525 2380 6325 2390
rect -70 2340 720 2350
rect -70 1170 -60 2340
rect 710 1170 720 2340
rect -70 1160 720 1170
rect 1530 2340 2320 2350
rect 1530 1170 1540 2340
rect 2310 1170 2320 2340
rect 1530 1160 2320 1170
rect 3130 2340 3920 2350
rect 3130 1170 3140 2340
rect 3910 1170 3920 2340
rect 3130 1160 3920 1170
rect 4730 2340 5520 2350
rect 4730 1170 4740 2340
rect 5510 1170 5520 2340
rect 4730 1160 5520 1170
rect 6330 2340 7120 2350
rect 6330 1170 6340 2340
rect 7110 1170 7120 2340
rect 6330 1160 7120 1170
rect 7930 2340 8720 3365
rect 9525 4535 10315 4545
rect 9525 3365 9535 4535
rect 10305 3365 10315 4535
rect 9525 3355 10315 3365
rect 10355 4535 11145 4545
rect 10355 3365 10365 4535
rect 11135 3365 11145 4535
rect 10355 3355 11145 3365
rect 11955 4535 12745 4545
rect 11955 3365 11965 4535
rect 12735 3365 12745 4535
rect 11955 3320 12745 3365
rect 13555 4535 14345 4770
rect 13555 3365 13565 4535
rect 14335 3365 14345 4535
rect 13555 3355 14345 3365
rect 11790 3255 12745 3320
rect 13590 3315 14345 3355
rect 13035 3280 14345 3315
rect 14385 5940 15175 5950
rect 14385 4770 14395 5940
rect 15165 4770 15175 5940
rect 14385 4535 15175 4770
rect 15985 5940 16775 5950
rect 15985 4770 15995 5940
rect 16765 4770 16775 5940
rect 15985 4760 16775 4770
rect 17585 5940 18375 5950
rect 17585 4770 17595 5940
rect 18365 4770 18375 5940
rect 17585 4760 18375 4770
rect 16780 4720 17580 4730
rect 16780 4700 16790 4720
rect 17570 4700 17580 4720
rect 16780 4690 17580 4700
rect 16780 4605 17580 4615
rect 16780 4585 16790 4605
rect 17570 4585 17580 4605
rect 16780 4575 17580 4585
rect 14385 3365 14395 4535
rect 15165 3365 15175 4535
rect 14385 3355 15175 3365
rect 15985 4535 16775 4545
rect 15985 3365 15995 4535
rect 16765 3365 16775 4535
rect 15985 3355 16775 3365
rect 17585 4535 18375 4545
rect 17585 3365 17595 4535
rect 18365 3365 18375 4535
rect 17585 3355 18375 3365
rect 9070 3240 10260 3250
rect 9070 2520 9080 3240
rect 10250 2520 10260 3240
rect 9070 2510 10260 2520
rect 11790 2510 11860 3255
rect 11790 2470 11805 2510
rect 11845 2470 11860 2510
rect 10325 2410 11125 2420
rect 10325 2390 10335 2410
rect 11115 2390 11125 2410
rect 11790 2400 11860 2470
rect 13035 2420 13075 3280
rect 13115 3250 14305 3260
rect 13115 2530 13125 3250
rect 14295 2530 14305 3250
rect 14385 3230 15140 3355
rect 14325 3220 15140 3230
rect 14325 3200 14345 3220
rect 15125 3200 15140 3220
rect 14325 3190 15140 3200
rect 16030 3260 16780 3355
rect 13115 2520 14305 2530
rect 16030 2460 16100 3260
rect 16280 3225 17470 3235
rect 16280 2505 16290 3225
rect 17460 2505 17470 3225
rect 16280 2495 17470 2505
rect 10325 2380 11125 2390
rect 11185 2350 11860 2400
rect 11925 2410 13075 2420
rect 11925 2390 11935 2410
rect 12715 2390 13075 2410
rect 11925 2380 13075 2390
rect 14860 2400 16100 2460
rect 14860 2350 15120 2400
rect 7930 1170 7940 2340
rect 8710 1170 8720 2340
rect 7930 1160 8720 1170
rect 9530 2340 10320 2350
rect 9530 1170 9540 2340
rect 10310 1170 10320 2340
rect 9530 1160 10320 1170
rect 11130 2340 11920 2350
rect 11130 1170 11140 2340
rect 11910 1170 11920 2340
rect 11130 1160 11920 1170
rect 12730 2340 13520 2350
rect 12730 1170 12740 2340
rect 13510 1170 13520 2340
rect 12730 1160 13520 1170
rect 14330 2340 15120 2350
rect 14330 1170 14340 2340
rect 15110 1170 15120 2340
rect 14330 1160 15120 1170
rect 15930 2340 16720 2350
rect 15930 1170 15940 2340
rect 16710 1170 16720 2340
rect 15930 1160 16720 1170
rect 725 1120 1525 1130
rect 725 1100 735 1120
rect 1515 1100 1525 1120
rect 725 1090 1525 1100
rect 1600 1110 2320 1160
rect 14330 1110 15050 1160
rect 1600 1065 15050 1110
rect 15125 1120 15925 1130
rect 15125 1100 15135 1120
rect 15915 1100 15925 1120
rect 15125 1090 15925 1100
<< viali >>
rect 735 8185 1515 8205
rect 15135 8185 15915 8205
rect -60 6965 710 8135
rect 3140 6965 3910 8135
rect 6340 6965 7110 8135
rect -810 6080 360 6800
rect 5535 6895 6315 6915
rect 2355 6055 3525 6775
rect 6400 6065 7570 6785
rect -1715 4770 -945 5940
rect -920 4700 -140 4720
rect -920 4585 -140 4605
rect -1715 3365 -945 4535
rect -810 2505 360 3225
rect 5515 4770 6285 5940
rect 9540 6965 10310 8135
rect 12740 6965 13510 8135
rect 10335 6895 11115 6915
rect 15940 6965 16710 8135
rect 9080 6065 10250 6785
rect 13125 6055 14295 6775
rect 10365 4770 11135 5940
rect 16290 6080 17460 6800
rect 4710 4700 5490 4720
rect 11160 4700 11940 4720
rect 4710 4585 5490 4605
rect 11160 4585 11940 4605
rect 5515 3365 6285 4535
rect 2355 2530 3525 3250
rect 6400 2520 7570 3240
rect 5535 2390 6315 2410
rect -60 1170 710 2340
rect 3140 1170 3910 2340
rect 6340 1170 7110 2340
rect 10365 3365 11135 4535
rect 17595 4770 18365 5940
rect 16790 4700 17570 4720
rect 16790 4585 17570 4605
rect 17595 3365 18365 4535
rect 9080 2520 10250 3240
rect 10335 2390 11115 2410
rect 13125 2530 14295 3250
rect 16290 2505 17460 3225
rect 9540 1170 10310 2340
rect 12740 1170 13510 2340
rect 15940 1170 16710 2340
rect 735 1100 1515 1120
rect 15135 1100 15915 1120
<< metal1 >>
rect -1790 8205 18445 8265
rect -1790 8185 735 8205
rect 1515 8185 15135 8205
rect 15915 8185 18445 8205
rect -1790 8135 18445 8185
rect -1790 6965 -60 8135
rect 710 6965 3140 8135
rect 3910 6965 6340 8135
rect 7110 6965 9540 8135
rect 10310 6965 12740 8135
rect 13510 6965 15940 8135
rect 16710 6965 18445 8135
rect -1790 6915 18445 6965
rect -1790 6895 5535 6915
rect 6315 6895 10335 6915
rect 11115 6895 18445 6915
rect -1790 6800 18445 6895
rect -1790 6080 -810 6800
rect 360 6785 16290 6800
rect 360 6775 6400 6785
rect 360 6080 2355 6775
rect -1790 6055 2355 6080
rect 3525 6065 6400 6775
rect 7570 6065 9080 6785
rect 10250 6775 16290 6785
rect 10250 6065 13125 6775
rect 3525 6055 13125 6065
rect 14295 6080 16290 6775
rect 17460 6080 18445 6800
rect 14295 6055 18445 6080
rect -1790 5940 18445 6055
rect -1790 4770 -1715 5940
rect -945 4770 5515 5940
rect 6285 4770 10365 5940
rect 11135 4770 17595 5940
rect 18365 4770 18445 5940
rect -1790 4720 18445 4770
rect -1790 4700 -920 4720
rect -140 4700 4710 4720
rect 5490 4700 11160 4720
rect 11940 4700 16790 4720
rect 17570 4700 18445 4720
rect -1790 4690 18445 4700
rect -1790 4605 18445 4620
rect -1790 4585 -920 4605
rect -140 4585 4710 4605
rect 5490 4585 11160 4605
rect 11940 4585 16790 4605
rect 17570 4585 18445 4605
rect -1790 4535 18445 4585
rect -1790 3365 -1715 4535
rect -945 3365 5515 4535
rect 6285 3365 10365 4535
rect 11135 3365 17595 4535
rect 18365 3365 18445 4535
rect -1790 3250 18445 3365
rect -1790 3225 2355 3250
rect -1790 2505 -810 3225
rect 360 2530 2355 3225
rect 3525 3240 13125 3250
rect 3525 2530 6400 3240
rect 360 2520 6400 2530
rect 7570 2520 9080 3240
rect 10250 2530 13125 3240
rect 14295 3225 18445 3250
rect 14295 2530 16290 3225
rect 10250 2520 16290 2530
rect 360 2505 16290 2520
rect 17460 2505 18445 3225
rect -1790 2410 18445 2505
rect -1790 2390 5535 2410
rect 6315 2390 10335 2410
rect 11115 2390 18445 2410
rect -1790 2340 18445 2390
rect -1790 1170 -60 2340
rect 710 1170 3140 2340
rect 3910 1170 6340 2340
rect 7110 1170 9540 2340
rect 10310 1170 12740 2340
rect 13510 1170 15940 2340
rect 16710 1170 18445 2340
rect -1790 1120 18445 1170
rect -1790 1100 735 1120
rect 1515 1100 15135 1120
rect 15915 1100 18445 1120
rect -1790 1080 18445 1100
<< labels >>
rlabel locali -1790 3285 -1790 3285 7 Idump
port 3 w
rlabel poly -1790 3150 -1790 3150 7 Vcn
port 4 w
rlabel poly -1790 2435 -1790 2435 7 Iout
port 5 w
rlabel poly -1790 6880 -1790 6880 7 Vbp
port 1 w
rlabel poly -1790 6020 -1790 6020 7 Vcp
port 2 w
rlabel metal1 -1790 6425 -1790 6425 7 VP
port 7 w
rlabel poly 18445 4655 18445 4655 3 Ifout
port 6 e
rlabel metal1 -1790 2811 -1790 2811 7 VN
<< end >>
