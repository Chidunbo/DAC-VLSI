* NGSPICE file created from cascode_voltage_gen.ext - technology: sky130A

X0 a_3140_3350# a_1540_3320# VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X1 a_3140_3350# a_1540_3320# VP VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X2 VP Vbp a_0_n30# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X3 VP Vbp Vcn VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=48 ps=28 w=6 l=8
X4 a_3140_3350# a_1540_3320# a_1540_3320# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X5 a_0_n30# a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X6 a_1600_0# Vcn Vcn VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X7 a_1600_0# Vcn Vcn VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X8 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=624 ps=364 w=6 l=8
X9 VP Vbp Vcn VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=48 ps=28 w=6 l=8
X10 a_1600_0# a_0_n30# VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X11 Vcp Vcp a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X12 a_1600_0# a_0_n30# a_0_n30# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X13 a_1540_3320# a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X14 a_1600_0# a_0_n30# a_0_n30# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X15 VN Vbn a_1540_3320# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X16 Vcn Vcn a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X17 a_3140_3350# Vcp Vcp VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X18 VP a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X19 VN a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X20 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=528 ps=308 w=6 l=8
X21 VP a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X22 a_1540_3320# a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X23 Vcp Vbn VN VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X24 a_3140_3350# Vcp Vcp VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X25 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=0 ps=0 w=6 l=8
X26 a_0_n30# a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X27 a_1600_0# a_0_n30# a_0_n30# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X28 VN a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X29 Vcp Vbn VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X30 a_1540_3320# a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X31 VN Vbn Vcp VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=48 ps=28 w=6 l=8
X32 VN Vbn Vcp VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X33 VN VN VN VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=0 ps=0 w=6 l=8
X34 a_3140_3350# a_1540_3320# a_1540_3320# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X35 a_1540_3320# a_1540_3320# a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X36 VN VN Vcp VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X37 a_0_n30# a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X38 a_0_n30# a_0_n30# a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X39 a_1600_0# a_0_n30# a_0_n30# VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X40 a_1540_3320# Vbn VN VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X41 Vcn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X42 Vcn Vbp VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=48 ps=28 w=6 l=8
X43 Vcn Vcn a_1600_0# VN sky130_fd_pr__nfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X44 a_0_n30# Vbp VP VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X45 Vcp Vcp a_3140_3350# VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=24 ps=14 w=6 l=8
X46 a_3140_3350# a_1540_3320# a_1540_3320# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=24 ps=14 w=6 l=8
X47 VP VP VP VP sky130_fd_pr__pfet_01v8 ad=48 pd=28 as=0 ps=0 w=6 l=8
X48 a_1600_0# a_0_n30# VN VN sky130_fd_pr__nfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8
X49 a_3140_3350# a_1540_3320# a_1540_3320# VP sky130_fd_pr__pfet_01v8 ad=24 pd=14 as=48 ps=28 w=6 l=8

